library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017
-- Dudy Nov 13 2017


entity back_ground_draw_new is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end back_ground_draw_new;

architecture behav of back_ground_draw_new is 

constant object_X_size : integer := 640;
constant object_Y_size : integer := 480;


type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  

constant object_colors: ram_array := ( 


     (x"ff",x"db",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b2",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"45",x"6d",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"8d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"6d",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"45",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"25",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"24",x"25",x"49",x"69",x"6d",x"6e",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"b2",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"b6",x"49",x"25",x"24",x"24",x"24",x"25",x"25",x"49",x"b6",x"b6",x"49",x"45",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"d7",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"fb",x"8d",x"69",x"69",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"d6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"db",x"db",x"db",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"b7",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"20",x"24",x"20",x"00",x"24",x"49",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"6d",x"69",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b6",x"b2",x"6d",x"69",x"49",x"49",x"69",x"6d",x"b2",x"db",x"db",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"45",x"25",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"45",x"45",x"6d",x"b6",x"6d",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b2",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"92",x"69",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"ff",x"fb",x"ff",x"db",x"ff",x"ff",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"25",x"49",x"db",x"b7",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"d7",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"8e",x"b6",x"92",x"49",x"24",x"45",x"25",x"24",x"25",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"49",x"6d",x"49",x"49",x"45",x"49",x"45",x"49",x"49",x"69",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"45",x"25",x"25",x"25",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"49",x"6d",x"b2",x"b6",x"92",x"92",x"92",x"92",x"b6",x"b6",x"db",x"db",x"b6",x"6d",x"49",x"45",x"45",x"45",x"45",x"45",x"49",x"49",x"24",x"45",x"49",x"92",x"6d",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"8e",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6e",x"6d",x"6e",x"92",x"b6",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"da",x"b6",x"b6",x"b6",x"b6",x"ff",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"69",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"fb",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"b6",x"b6",x"ff",x"b6",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"25",x"24",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"b7",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"49",x"49",x"45",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"25",x"24",x"25",x"45",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"92",x"b6",x"d7",x"b6",x"d6",x"b6",x"b6",x"b2",x"92",x"b2",x"b7",x"92",x"49",x"24",x"24",x"25",x"45",x"45",x"24",x"45",x"45",x"49",x"49",x"92",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"6e",x"6d",x"6d",x"6d",x"6e",x"b2",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"da",x"b6",x"b6",x"b6",x"da",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"6d",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"8d",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"49",x"49",x"24",x"24",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"b6",x"fb",x"b6",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"25",x"6d",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"8e",x"49",x"49",x"45",x"25",x"45",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"92",x"d7",x"d7",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"45",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"b6",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"92",x"db",x"92",x"6d",x"49",x"49",x"69",x"6d",x"92",x"b6",x"ff",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"da",x"b6",x"b6",x"d6",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"6d",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"8e",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"92",x"92",x"92",x"8e",x"92",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"49",x"92",x"db",x"92",x"92",x"92",x"92",x"b6",x"db",x"fb",x"db",x"b2",x"49",x"49",x"49",x"45",x"44",x"25",x"25",x"24",x"25",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6e",x"6e",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"69",x"49",x"45",x"45",x"49",x"49",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"49",x"49",x"45",x"45",x"49",x"6d",x"b6",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"da",x"b6",x"b6",x"da",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"69",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"6d",x"8d",x"92",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"8e",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"d7",x"6d",x"69",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"b6",x"d7",x"8e",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"25",x"45",x"24",x"24",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"20",x"20",x"45",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"69",x"49",x"6d",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"8e",x"b2",x"6d",x"49",x"45",x"45",x"25",x"25",x"25",x"49",x"8e",x"92",x"69",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"92",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"da",x"b6",x"b6",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"8d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"49",x"49",x"6d",x"da",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"b2",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"6d",x"69",x"49",x"49",x"69",x"6d",x"92",x"b6",x"8d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"25",x"24",x"45",x"24",x"45",x"49",x"24",x"24",x"6d",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"6e",x"92",x"6d",x"49",x"49",x"49",x"49",x"6e",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"92",x"92",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"8e",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"8e",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"25",x"25",x"25",x"45",x"45",x"25",x"45",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"8d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"da",x"db",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b2",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"69",x"b2",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"6d",x"6e",x"49",x"49",x"49",x"49",x"25",x"45",x"45",x"49",x"6d",x"6d",x"49",x"49",x"45",x"45",x"45",x"24",x"25",x"25",x"25",x"24",x"24",x"6d",x"b2",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"6d",x"6e",x"49",x"24",x"24",x"49",x"6d",x"92",x"92",x"b2",x"b2",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6e",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"45",x"25",x"49",x"49",x"6d",x"49",x"49",x"45",x"49",x"6d",x"6d",x"49",x"49",x"45",x"44",x"44",x"49",x"6d",x"92",x"6e",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"25",x"24",x"24",x"25",x"24",x"25",x"45",x"25",x"45",x"45",x"49",x"6d",x"92",x"49",x"24",x"45",x"45",x"45",x"49",x"45",x"45",x"49",x"92",x"b7",x"92",x"69",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"69",x"49",x"69",x"6d",x"6d",x"92",x"b6",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"db",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ba",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"b6",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"69",x"b2",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"49",x"49",x"45",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"92",x"b7",x"92",x"69",x"45",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"25",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"45",x"20",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"92",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"92",x"6d",x"6d",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"45",x"45",x"49",x"49",x"6d",x"6d",x"24",x"24",x"45",x"45",x"45",x"45",x"24",x"45",x"45",x"49",x"b6",x"b6",x"92",x"6d",x"69",x"6d",x"6d",x"92",x"db",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"db",x"b6",x"db",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"69",x"49",x"6d",x"6d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b2",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"25",x"45",x"49",x"45",x"25",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"b6",x"b2",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"20",x"24",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"45",x"25",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"6d",x"8e",x"8e",x"8e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"b2",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"69",x"49",x"24",x"24",x"49",x"6d",x"b2",x"b6",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"45",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"45",x"49",x"49",x"92",x"d7",x"d7",x"b6",x"92",x"92",x"b6",x"db",x"fb",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"fb",x"db",x"fb",x"ff",x"ff",x"ff",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"fb",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b2",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"da",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"fb",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"d6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6e",x"49",x"49",x"49",x"25",x"45",x"49",x"45",x"25",x"24",x"49",x"6d",x"49",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"6d",x"8e",x"92",x"92",x"92",x"b6",x"b6",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"69",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"20",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"92",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"25",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"6d",x"69",x"49",x"24",x"24",x"25",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"92",x"6d",x"6d",x"6d",x"8e",x"92",x"92",x"6e",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"25",x"25",x"24",x"49",x"49",x"45",x"45",x"49",x"49",x"6d",x"d7",x"db",x"db",x"db",x"b7",x"db",x"db",x"db",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6"),
     (x"49",x"49",x"49",x"49",x"d6",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"db",x"db",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"d7",x"6d",x"49",x"49",x"49",x"49",x"45",x"25",x"25",x"45",x"24",x"49",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"6e",x"6d",x"49",x"25",x"49",x"49",x"6d",x"b2",x"b6",x"b2",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"8e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b2",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"24",x"24",x"24",x"25",x"49",x"45",x"45",x"49",x"92",x"49",x"25",x"45",x"25",x"45",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"b6",x"db",x"db",x"d7",x"b6",x"b6",x"b2",x"b6",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"ff",x"db",x"b6",x"92",x"b2",x"b2",x"b6",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"91",x"b6",x"d6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"ff",x"92",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"d6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"8e",x"6d",x"6d",x"6d",x"b2",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"24",x"45",x"92",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"6e",x"6d",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"45",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"25",x"49",x"24",x"20",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"49",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"6d",x"92",x"6e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"6d",x"b6",x"49",x"24",x"45",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"8e",x"6d",x"6d",x"6d",x"8e",x"b6",x"d7",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"db",x"b6",x"8e",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"92",x"db",x"b6",x"6d",x"69",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"6d",x"fb",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"d6",x"b2",x"92",x"8d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"45",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"b6",x"b2",x"b6",x"b6",x"db",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"45",x"8e",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"45",x"6d",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"20",x"20",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"45",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"92",x"49",x"45",x"24",x"24",x"45",x"49",x"6d",x"b6",x"b6",x"69",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"d7",x"8e",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"fb",x"b6",x"92",x"91",x"92",x"92",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"db",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"8e",x"92",x"b6",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"69",x"db",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"b6",x"8e",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"db",x"6d",x"49",x"49",x"45",x"49",x"24",x"45",x"49",x"25",x"49",x"45",x"49",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"45",x"49",x"92",x"b6",x"8e",x"49",x"49",x"45",x"45",x"45",x"49",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"24",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"25",x"24",x"49",x"49",x"69",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b7",x"b6",x"6d",x"25",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"b2",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"fb",x"db",x"b2",x"92",x"92",x"b2",x"b6",x"ff",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"92",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"ff",x"d7",x"92",x"92",x"92",x"b6",x"db",x"ff",x"fb",x"6d",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"24",x"49",x"25",x"49",x"db",x"fb",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"45",x"24",x"25",x"92",x"db",x"b6",x"92",x"69",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"69",x"25",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"04",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"20",x"24",x"24",x"20",x"24",x"20",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"45",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"b6",x"b6",x"6d",x"45",x"45",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"92",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"44",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"db",x"b6",x"b6",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"db",x"b6",x"b6",x"db",x"ff",x"ff",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"25",x"49",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"45",x"24",x"24",x"92",x"d7",x"d7",x"b6",x"b2",x"92",x"b2",x"b6",x"d7",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b7",x"b6",x"b6",x"92",x"6e",x"6d",x"6e",x"b2",x"92",x"49",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"b2",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"fb",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"24",x"24",x"45",x"45",x"45",x"45",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"92",x"92",x"8e",x"6d",x"92",x"92",x"b6",x"d7",x"b6",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6e",x"8e",x"69",x"45",x"24",x"24",x"45",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"00",x"24",x"25",x"45",x"25",x"25",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"92",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"92",x"6e",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"69",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"45",x"49",x"49",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"92",x"92",x"69",x"49",x"45",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"db",x"ff",x"ff",x"fb",x"fb",x"db",x"fb",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"d6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"ff",x"db",x"db",x"b7",x"db",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"4d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"db",x"d6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"8e",x"49",x"24",x"24",x"44",x"24",x"24",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"db",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"49",x"69",x"6e",x"8e",x"6d",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"00",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"20",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"69",x"6d",x"49",x"45",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"45",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"8e",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"92",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"db",x"b7",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"6d",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"24",x"24",x"44",x"44",x"49",x"49",x"49",x"49",x"6d",x"fb",x"ff",x"db",x"db",x"b6",x"b6",x"b2",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"00",x"00",x"49",x"6d",x"69",x"49",x"49",x"49",x"45",x"24",x"24",x"25",x"20",x"00",x"00",x"24",x"24",x"20",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"92",x"92",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"92",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"20",x"00",x"20",x"20",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"45",x"45",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"44",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"b2",x"ff",x"db",x"b6",x"b6",x"d7",x"db",x"ff",x"ff",x"ff",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"45",x"b6",x"92",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"fb",x"fb",x"ff",x"db",x"db",x"ff",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"25",x"24",x"44",x"24",x"25",x"49",x"49",x"49",x"49",x"db",x"ff",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"b2",x"db",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"69",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"8e",x"49",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"20",x"20",x"20",x"24",x"49",x"45",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"8e",x"49",x"49",x"49",x"49",x"45",x"25",x"45",x"49",x"49",x"49",x"b2",x"db",x"92",x"69",x"49",x"49",x"49",x"6d",x"8e",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"d7",x"db",x"b6",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"ff",x"db",x"db",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"24",x"92",x"b6",x"49",x"49",x"44",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"da",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"db",x"ff",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"69",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"92",x"92",x"6d",x"49",x"49",x"69",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"20",x"20",x"00",x"00",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"8e",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"20",x"20",x"24",x"25",x"24",x"00",x"00",x"00",x"20",x"20",x"00",x"20",x"24",x"20",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"00",x"20",x"20",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"8e",x"69",x"49",x"25",x"49",x"49",x"6e",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"49",x"49",x"92",x"db",x"d7",x"8d",x"6d",x"6d",x"6d",x"8d",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"8e",x"db",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"69",x"b6",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"96",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"fb",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"db",x"6e",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"45",x"45",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"92",x"b2",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"25",x"25",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"24",x"20",x"20",x"20",x"20",x"24",x"24",x"20",x"00",x"20",x"20",x"00",x"20",x"24",x"24",x"20",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"92",x"92",x"6e",x"6d",x"69",x"49",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b6",x"b6",x"6d",x"49",x"69",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"fb",x"b6",x"92",x"8d",x"92",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"6d",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"92",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"b6",x"6d",x"49",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"fb",x"db",x"b6",x"92",x"b6",x"db",x"db",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"45",x"49",x"25",x"45",x"45",x"49",x"49",x"49",x"45",x"8e",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"25",x"24",x"20",x"00",x"20",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"20",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"25",x"25",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"6d",x"49",x"25",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"45",x"69",x"b6",x"d7",x"b6",x"92",x"92",x"b6",x"db",x"db",x"b6",x"69",x"45",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"d7",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"25",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"96",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"6d",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"92",x"92",x"49",x"44",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"24",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ba",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"b2",x"db",x"6d",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"45",x"49",x"45",x"49",x"49",x"49",x"45",x"69",x"d7",x"92",x"69",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"49",x"25",x"24",x"24",x"20",x"24",x"20",x"20",x"20",x"24",x"49",x"24",x"20",x"24",x"20",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"8e",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"45",x"49",x"b2",x"d7",x"d7",x"b6",x"b6",x"b6",x"d7",x"db",x"b7",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"db",x"db",x"db",x"db",x"fb",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"45",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"69",x"69",x"49",x"6d",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"b6",x"8d",x"6d",x"6d",x"92",x"92",x"92",x"db",x"ff",x"db",x"b6",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"6d",x"b6",x"49",x"44",x"24",x"49",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"d6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"b6",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"45",x"45",x"45",x"25",x"49",x"45",x"49",x"d7",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"d7",x"b6",x"6d",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"49",x"69",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"45",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"45",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"25",x"49",x"25",x"25",x"45",x"45",x"49",x"92",x"b6",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"d7",x"69",x"45",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"db",x"b6",x"b6",x"b6",x"d7",x"db",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"6d",x"69",x"49",x"49",x"49",x"69",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"db",x"92",x"92",x"91",x"91",x"92",x"92",x"b6",x"db",x"db",x"b6",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"92",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"b6",x"6d",x"48",x"24",x"49",x"24",x"49",x"49",x"48",x"24",x"24",x"24",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"df",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"91",x"b6",x"d6",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"49",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"45",x"49",x"45",x"45",x"b2",x"ff",x"db",x"b6",x"b2",x"b6",x"d7",x"db",x"d7",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"49",x"69",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"49",x"69",x"6d",x"49",x"49",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"92",x"6e",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"44",x"24",x"44",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"49",x"49",x"69",x"8e",x"92",x"8e",x"45",x"24",x"24",x"24",x"25",x"49",x"45",x"45",x"45",x"45",x"69",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"b6",x"92",x"6e",x"8e",x"92",x"92",x"db",x"db",x"92",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"49",x"49",x"49",x"92",x"fb",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"b2",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"49",x"49",x"49",x"45",x"45",x"49",x"45",x"49",x"49",x"49",x"69",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"48",x"24",x"24",x"24",x"49",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"92",x"8e",x"6d",x"6d",x"6d",x"92",x"d6",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"45",x"24",x"24",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"b6",x"fb",x"6e",x"49",x"49",x"49",x"49",x"45",x"24",x"25",x"24",x"25",x"45",x"92",x"db",x"db",x"b6",x"b6",x"b6",x"d7",x"db",x"b6",x"49",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"20",x"20",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"25",x"24",x"45",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"6d",x"b2",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"b2",x"92",x"8e",x"8e",x"92",x"92",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"25",x"45",x"45",x"45",x"6d",x"6e",x"49",x"49",x"45",x"25",x"25",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"b6",x"6e",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"d6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"92",x"db",x"ff",x"db",x"96",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"d6",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"6d",x"69",x"6d",x"92",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"45",x"24",x"8e",x"b6",x"92",x"8e",x"6d",x"6e",x"8e",x"92",x"92",x"69",x"25",x"45",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"92",x"92",x"92",x"92",x"b6",x"b6",x"8e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"6d",x"69",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"45",x"25",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"24",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6e",x"92",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"69",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"49",x"25",x"25",x"25",x"25",x"25",x"45",x"49",x"92",x"6d",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"45",x"24",x"45",x"25",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"24",x"49",x"44",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"48",x"24",x"24",x"24",x"49",x"49",x"45",x"44",x"24",x"24",x"6e",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"d6",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"8d",x"da",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"b6",x"92",x"8d",x"92",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"45",x"49",x"49",x"45",x"24",x"45",x"24",x"24",x"24",x"24",x"8e",x"6d",x"49",x"49",x"6d",x"6e",x"92",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6e",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"25",x"24",x"49",x"6d",x"6d",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"45",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"20",x"00",x"20",x"00",x"20",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"20",x"20",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"6d",x"49",x"24",x"00",x"20",x"20",x"20",x"20",x"24",x"45",x"49",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"45",x"25",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"6e",x"6d",x"45",x"24",x"24",x"25",x"25",x"45",x"49",x"49",x"49",x"6d",x"49",x"25",x"25",x"25",x"25",x"45",x"45",x"49",x"92",x"92",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"fb",x"b2",x"91",x"6d",x"8d",x"92",x"b6",x"db",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"49",x"49",x"49",x"45",x"44",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b2",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"db",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"b6",x"6d",x"49",x"24",x"44",x"24",x"44",x"49",x"45",x"49",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"b6",x"db",x"b2",x"92",x"8d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"d6",x"b6",x"b6",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"45",x"24",x"6d",x"8e",x"49",x"25",x"45",x"25",x"44",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"25",x"49",x"24",x"24",x"25",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"25",x"25",x"24",x"24",x"45",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"24",x"00",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"6d",x"6d",x"49",x"25",x"24",x"25",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"45",x"49",x"45",x"25",x"45",x"45",x"6d",x"49",x"25",x"25",x"25",x"24",x"25",x"45",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"6d",x"49",x"69",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff"),
     (x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"d6",x"92",x"92",x"92",x"92",x"b2",x"db",x"ff",x"ff",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"45",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"25",x"25",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"6d",x"49",x"24",x"25",x"24",x"45",x"25",x"24",x"49",x"6d",x"6e",x"92",x"6d",x"49",x"24",x"49",x"45",x"25",x"25",x"25",x"24",x"49",x"49",x"45",x"25",x"49",x"24",x"25",x"49",x"24",x"49",x"49",x"25",x"25",x"49",x"49",x"25",x"49",x"49",x"25",x"45",x"45",x"45",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"45",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"45",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"49",x"24",x"25",x"25",x"24",x"24",x"25",x"45",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db"),
     (x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"48",x"24",x"44",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"db",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"45",x"45",x"49",x"db",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"25",x"45",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"8e",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"69",x"8e",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"6d",x"6d",x"25",x"24",x"25",x"25",x"24",x"25",x"25",x"25",x"49",x"92",x"92",x"92",x"92",x"92",x"b6",x"92",x"49",x"24",x"45",x"24",x"25",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"20",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"49",x"49",x"45",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"49",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"69",x"6d",x"49",x"25",x"45",x"25",x"24",x"24",x"25",x"25",x"45",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"8e"),
     (x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"6d",x"49",x"44",x"44",x"24",x"45",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"db",x"b6",x"b2",x"b6",x"db",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"49",x"24",x"45",x"25",x"24",x"49",x"6d",x"49",x"45",x"45",x"49",x"49",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"6d",x"8e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"25",x"25",x"25",x"25",x"25",x"25",x"25",x"6d",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"25",x"49",x"25",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"69",x"49",x"24",x"24",x"25",x"49",x"25",x"49",x"49",x"92",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"8e",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"92",x"49",x"49",x"45",x"49",x"49",x"69",x"92",x"6d",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"25",x"25",x"6d",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6d",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"db",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d"),
     (x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"92",x"92",x"49",x"48",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"49",x"49",x"49",x"b6",x"db",x"92",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"db",x"b6",x"8e",x"6d",x"49",x"49",x"49",x"6e",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"6e",x"49",x"45",x"49",x"25",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"25",x"25",x"24",x"24",x"49",x"69",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"49",x"45",x"24",x"24",x"49",x"6d",x"49",x"49",x"45",x"24",x"24",x"25",x"49",x"6d",x"49",x"6d",x"6d",x"6e",x"8e",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"49",x"45",x"49",x"92",x"49",x"24",x"49",x"25",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"69",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"45",x"6d",x"d7",x"b6",x"6d",x"69",x"49",x"69",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"25",x"25",x"6d",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"db",x"b6",x"b6",x"db",x"fb",x"ff",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"45",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b2",x"b6",x"db",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49"),
     (x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"48",x"44",x"45",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"6e",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"fb",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"8e",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"49",x"24",x"24",x"24",x"25",x"45",x"25",x"49",x"92",x"6d",x"49",x"45",x"45",x"45",x"49",x"6d",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"25",x"24",x"49",x"69",x"49",x"25",x"24",x"00",x"00",x"00",x"24",x"49",x"6d",x"49",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"6e",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"25",x"69",x"8e",x"6d",x"6d",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"25",x"25",x"49",x"49",x"25",x"25",x"24",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"24",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"25",x"25",x"24",x"24",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"92",x"b6",x"92",x"92",x"92",x"b2",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"6d",x"b7",x"db",x"b2",x"8d",x"6d",x"8d",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"25",x"45",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"b7",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49"),
     (x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"b6",x"6d",x"49",x"48",x"49",x"24",x"48",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"fb",x"db",x"db",x"b6",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"8d",x"b6",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"45",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"00",x"20",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"25",x"25",x"25",x"49",x"49",x"49",x"92",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"49",x"6d",x"6d",x"69",x"49",x"25",x"24",x"49",x"49",x"45",x"49",x"49",x"6e",x"b6",x"6d",x"49",x"25",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"6d",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"92",x"b2",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"25",x"25",x"49",x"49",x"6e",x"d7",x"db",x"d7",x"b6",x"b2",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"25",x"45",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"db",x"b6",x"8e",x"6d",x"8e",x"92",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"92",x"92",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69"),
     (x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"8d",x"db",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"25",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"6e",x"b7",x"b6",x"92",x"8e",x"92",x"b2",x"db",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"8e",x"49",x"45",x"45",x"45",x"49",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"b2",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"25",x"24",x"49",x"25",x"25",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"b6",x"6e",x"25",x"25",x"25",x"45",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"45",x"49",x"49",x"45",x"25",x"24",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"45",x"25",x"25",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6e",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"69",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"45",x"49",x"49",x"92",x"b7",x"d7",x"d7",x"d7",x"d7",x"db",x"db",x"d7",x"69",x"49",x"49",x"45",x"25",x"45",x"49",x"45",x"25",x"45",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"d7",x"8e",x"6d",x"6d",x"6d",x"8e",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"45",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"92",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"db",x"b6",x"b6",x"d6",x"db",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d"),
     (x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"db",x"b2",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"8e",x"db",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"db",x"d7",x"b6",x"b6",x"b6",x"b6",x"b6",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"92",x"8e",x"6d",x"6e",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"25",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6e",x"6d",x"6d",x"6d",x"6d",x"69",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"45",x"45",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"20",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"49",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"49",x"49",x"25",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"92",x"6e",x"6d",x"6e",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"b2",x"b2",x"92",x"92",x"92",x"b2",x"b7",x"db",x"b6",x"49",x"49",x"49",x"25",x"25",x"25",x"25",x"25",x"24",x"49",x"92",x"db",x"6d",x"49",x"49",x"69",x"69",x"6d",x"6d",x"6d",x"d6",x"92",x"6d",x"6d",x"69",x"6d",x"6d",x"92",x"db",x"ff",x"6e",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"24",x"24",x"49",x"b6",x"6d",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"8d",x"91",x"92",x"b6",x"ff",x"ff",x"db",x"db",x"ff",x"db",x"db",x"b6",x"b6",x"db",x"ff",x"db",x"b6",x"92",x"92",x"6d",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d"),
     (x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b2",x"db",x"6e",x"45",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6e",x"6d",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"6d",x"8e",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"20",x"24",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"25",x"24",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"92",x"92",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"69",x"69",x"6d",x"92",x"b7",x"b2",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"25",x"25",x"49",x"b6",x"db",x"6d",x"69",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"69",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"db",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"db",x"da",x"db",x"db",x"ff",x"db",x"92",x"92",x"8d",x"6d",x"6d",x"92",x"d7",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"49",x"45",x"45",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"8e",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"6d",x"49",x"45",x"25",x"45",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"24",x"20",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"69",x"92",x"49",x"49",x"49",x"24",x"25",x"49",x"6d",x"92",x"6d",x"49",x"25",x"25",x"49",x"49",x"49",x"92",x"b2",x"6e",x"6e",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"45",x"49",x"25",x"24",x"49",x"6d",x"6e",x"92",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"29",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"20",x"20",x"20",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"25",x"49",x"25",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"d6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"44",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"91",x"92",x"92",x"b2",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"db",x"b6",x"92",x"8e",x"6d",x"6d",x"6d",x"b2",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"ff",x"b6",x"8e",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"44",x"44",x"25",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"b2",x"b2",x"b7",x"db",x"db",x"92",x"49",x"49",x"45",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"25",x"45",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"20",x"00",x"25",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"49",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"4d",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"25",x"49",x"49",x"49",x"6d",x"92",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"6d",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"49",x"49",x"69",x"db",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"ff",x"da",x"92",x"6d",x"6d",x"8d",x"92",x"92",x"92",x"d6",x"ff",x"db",x"b7",x"b7",x"db",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"92",x"ff",x"fb",x"db",x"db",x"db",x"db",x"b6",x"92",x"49",x"49",x"49",x"45",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"20",x"20",x"24",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"25",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"69",x"24",x"24",x"24",x"24",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"25",x"25",x"25",x"49",x"45",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"b2",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"45",x"49",x"49",x"25",x"6d",x"6d",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"20",x"6d",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"45",x"24",x"44",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"b6",x"6d",x"25",x"24",x"25",x"25",x"24",x"25",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"92",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"44",x"24",x"24",x"49",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"db",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"92",x"92",x"92",x"b2",x"ff",x"db",x"db",x"b6",x"b7",x"db",x"ff",x"ff",x"db",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b7",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"92",x"8d",x"6d",x"92",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"25",x"69",x"db",x"ff",x"db",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"45",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"49",x"45",x"24",x"24",x"20",x"24",x"24",x"25",x"49",x"25",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"25",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"49",x"25",x"49",x"49",x"25",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"69",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"69",x"49",x"6d",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6e",x"25",x"24",x"24",x"24",x"25",x"49",x"25",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"25",x"24",x"24",x"20",x"20",x"00",x"00",x"20",x"20",x"24",x"24",x"04",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"49",x"49",x"45",x"25",x"49",x"92",x"49",x"24",x"24",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"b2",x"fb",x"ff",x"d7",x"92",x"92",x"92",x"92",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"25",x"24",x"24",x"44",x"44",x"45",x"24",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"91",x"91",x"91",x"92",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"b6",x"b7",x"db",x"ff",x"ff",x"db",x"fb",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"b6",x"8e",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"24",x"24",x"24",x"6e",x"b6",x"25",x"25",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"db",x"b6",x"b2",x"92",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"b6",x"db",x"b6",x"92",x"6d",x"49",x"49",x"69",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"24",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"20",x"24",x"25",x"49",x"69",x"69",x"25",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"45",x"25",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"92",x"92",x"b6",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"b6",x"b2",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"25",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"45",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"25",x"20",x"00",x"00",x"00",x"20",x"20",x"24",x"49",x"24",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"8e",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"92",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"49",x"49",x"49",x"45",x"45",x"25",x"49",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"fb",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"44",x"49",x"92",x"d6",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"b2",x"fb",x"db",x"b6",x"b6",x"b6",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"92",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"44",x"44",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"fb",x"d6",x"b6",x"b2",x"b6",x"db",x"ff",x"db",x"ff",x"db",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"92",x"24",x"24",x"25",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"69",x"49",x"49",x"49",x"49",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"8e",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"45",x"25",x"49",x"49",x"6d",x"92",x"49",x"45",x"24",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"25",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"25",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"6e",x"69",x"49",x"69",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"92",x"b6",x"6e",x"49",x"49",x"49",x"49",x"6e",x"92",x"49",x"45",x"49",x"45",x"25",x"25",x"25",x"24",x"49",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"91",x"db",x"ff",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"b6",x"b6",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"8e",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"44",x"44",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"25",x"25",x"45",x"49",x"25",x"45",x"49",x"24",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"db",x"db",x"b6",x"db",x"db",x"db",x"db",x"db",x"db",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"49",x"49",x"6e",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"25",x"25",x"49",x"6d",x"49",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"8e",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"45",x"49",x"49",x"25",x"25",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"b6",x"b6",x"b6",x"b6",x"6e",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"24",x"25",x"49",x"25",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"24",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"25",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"92",x"6e",x"92",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"45",x"92",x"d7",x"92",x"6d",x"69",x"6d",x"92",x"b6",x"6d",x"25",x"49",x"45",x"25",x"24",x"25",x"25",x"25",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"92",x"b6",x"d7",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"48",x"44",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"49",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"db",x"fb",x"db",x"db",x"b6",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"49",x"25",x"45",x"25",x"49",x"49",x"45",x"69",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"b6",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"8e",x"8e",x"92",x"b6",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"49",x"49",x"49",x"6e",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"24",x"24",x"49",x"6d",x"49",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"24",x"00",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"45",x"49",x"25",x"24",x"25",x"49",x"6d",x"25",x"25",x"49",x"49",x"45",x"25",x"6d",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"92",x"92",x"b6",x"b6",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"6d",x"45",x"25",x"24",x"24",x"24",x"24",x"49",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"49",x"49",x"49",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"92",x"b7",x"b6",x"b2",x"92",x"b6",x"b6",x"92",x"49",x"25",x"25",x"25",x"24",x"24",x"25",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"b7",x"92",x"6d",x"92",x"b6",x"db",x"fb",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"49",x"b6",x"49",x"45",x"49",x"45",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b2",x"d6",x"ff",x"b6",x"b2",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"ff",x"ff",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"48",x"48",x"24",x"24",x"24",x"24",x"6d",x"b6",x"25",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"b2",x"92",x"b6",x"b6",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"45",x"25",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"49",x"24",x"25",x"25",x"49",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"24",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"6d",x"6d",x"6e",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"25",x"24",x"24",x"25",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"92",x"92",x"b2",x"92",x"b6",x"b6",x"6e",x"25",x"25",x"24",x"24",x"24",x"25",x"45",x"49",x"25",x"6d",x"b2",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b2",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"b6",x"49",x"49",x"49",x"45",x"49",x"45",x"45",x"25",x"24",x"6d",x"92",x"25",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"ff",x"ff",x"ff",x"ff",x"da",x"b6",x"92",x"92",x"b2",x"b6",x"fb",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"48",x"48",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"48",x"44",x"24",x"44",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"8d",x"b6",x"b6",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"45",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"6d",x"49",x"24",x"25",x"25",x"45",x"49",x"45",x"25",x"69",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"20",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"25",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"49",x"6d",x"b6",x"b2",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"69",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"b2",x"69",x"49",x"25",x"49",x"49",x"6d",x"b6",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"25",x"24",x"00",x"00",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"45",x"45",x"92",x"b2",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"b6",x"fb",x"8e",x"49",x"49",x"49",x"25",x"49",x"25",x"25",x"24",x"24",x"92",x"92",x"24",x"49",x"44",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"b6",x"92",x"b2",x"b6",x"da",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"da",x"6d",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"48",x"48",x"24",x"44",x"24",x"24",x"92",x"8d",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"b2",x"fb",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"25",x"25",x"24",x"49",x"49",x"25",x"45",x"b2",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"db",x"8e",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"20",x"20",x"24",x"00",x"20",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"45",x"24",x"00",x"00",x"00",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"6e",x"6e",x"25",x"49",x"49",x"49",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"8e",x"6d",x"6e",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"69",x"49",x"49",x"69",x"49",x"49",x"92",x"b6",x"92",x"92",x"92",x"92",x"6e",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"b6",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"49",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"45",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"24",x"20",x"20",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"6d",x"49",x"25",x"25",x"45",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"44",x"45",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"49",x"45",x"49",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"b6",x"69",x"44",x"49",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"d6",x"b6",x"b6",x"b6",x"b6",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff"),
     (x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"48",x"49",x"24",x"44",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"6e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b2",x"b6",x"92",x"6d",x"6d",x"6d",x"69",x"69",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"49",x"25",x"45",x"49",x"49",x"24",x"69",x"db",x"b6",x"92",x"92",x"b6",x"d7",x"db",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"20",x"20",x"24",x"24",x"04",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"20",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"49",x"b6",x"25",x"25",x"25",x"49",x"49",x"24",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"25",x"29",x"49",x"49",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"b6",x"d7",x"6d",x"69",x"69",x"69",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"25",x"49",x"25",x"25",x"24",x"24",x"24",x"45",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"d6",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff"),
     (x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"48",x"49",x"49",x"24",x"49",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"44",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"8d",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"24",x"24",x"49",x"6e",x"24",x"49",x"49",x"45",x"24",x"45",x"45",x"24",x"49",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"b2",x"92",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"69",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"20",x"20",x"00",x"00",x"25",x"49",x"24",x"24",x"20",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"69",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"49",x"25",x"25",x"49",x"6d",x"25",x"25",x"25",x"49",x"24",x"49",x"49",x"49",x"25",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"69",x"92",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"45",x"49",x"49",x"6d",x"6d",x"49",x"49",x"24",x"25",x"25",x"49",x"69",x"25",x"49",x"25",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"20",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"d7",x"db",x"92",x"6d",x"69",x"6d",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6e",x"24",x"45",x"45",x"49",x"24",x"24",x"24",x"45",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"db",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"da",x"ff",x"db",x"92",x"92",x"6d",x"6e",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db"),
     (x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"48",x"48",x"49",x"44",x"49",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"b2",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"db",x"d7",x"b2",x"92",x"6d",x"69",x"6d",x"69",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"20",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"6d",x"49",x"45",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"92",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"00",x"24",x"20",x"24",x"24",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"6d",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"45",x"25",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"25",x"45",x"45",x"49",x"49",x"92",x"db",x"db",x"b2",x"6d",x"6d",x"6d",x"8e",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"24",x"45",x"45",x"49",x"45",x"24",x"24",x"49",x"49",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"91",x"92",x"b6",x"ff",x"db",x"db",x"db",x"ff",x"db",x"da",x"b6",x"db",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92"),
     (x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"48",x"48",x"49",x"49",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"45",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"d7",x"92",x"8d",x"6d",x"92",x"db",x"ff",x"ff",x"d7",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"b6",x"92",x"b6",x"92",x"49",x"6d",x"49",x"49",x"49",x"92",x"49",x"69",x"69",x"6d",x"49",x"92",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"24",x"6d",x"6d",x"92",x"6d",x"24",x"24",x"49",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"45",x"24",x"24",x"00",x"20",x"49",x"24",x"00",x"20",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"20",x"20",x"20",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"49",x"69",x"b6",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"6e",x"b6",x"24",x"24",x"49",x"45",x"25",x"49",x"24",x"24",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"8d",x"92",x"92",x"db",x"db",x"db",x"b7",x"db",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"6d"),
     (x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"44",x"92",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"b6",x"92",x"b6",x"db",x"db",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"45",x"45",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"49",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"6e",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"92",x"69",x"45",x"49",x"49",x"25",x"49",x"b6",x"49",x"49",x"25",x"49",x"49",x"25",x"72",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"b6",x"db",x"92",x"49",x"69",x"49",x"69",x"49",x"6d",x"db",x"92",x"92",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"24",x"25",x"24",x"45",x"49",x"49",x"92",x"24",x"49",x"24",x"49",x"45",x"49",x"92",x"24",x"24",x"24",x"24",x"45",x"49",x"45",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"20",x"20",x"24",x"20",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"6e",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"92",x"49",x"45",x"25",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"69",x"24",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"db",x"db",x"b6",x"b6",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"92",x"6e",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"d6",x"ff",x"ff",x"db",x"92",x"8d",x"8d",x"8e",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"b6",x"db",x"ff",x"db",x"db",x"db",x"fb",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d"),
     (x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"44",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"49",x"25",x"49",x"25",x"49",x"49",x"24",x"92",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"fb",x"db",x"db",x"db",x"db",x"db",x"b6",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"6d",x"6d",x"92",x"b2",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"25",x"b6",x"24",x"24",x"25",x"25",x"49",x"24",x"6d",x"49",x"24",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"6e",x"6d",x"49",x"49",x"49",x"69",x"6e",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"69",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"45",x"49",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"25",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"20",x"20",x"24",x"20",x"20",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"b6",x"92",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"92",x"69",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"d7",x"b2",x"b6",x"db",x"db",x"db",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"25",x"25",x"92",x"49",x"24",x"24",x"24",x"45",x"45",x"45",x"24",x"49",x"49",x"b2",x"b6",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"91",x"92",x"92",x"92",x"b2",x"fb",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49"),
     (x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"da",x"49",x"44",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"92",x"24",x"24",x"49",x"24",x"25",x"24",x"25",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"49",x"45",x"45",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"20",x"24",x"45",x"49",x"24",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"45",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"45",x"25",x"49",x"24",x"6d",x"24",x"25",x"25",x"25",x"49",x"69",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"49",x"db",x"db",x"b6",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"b6",x"db",x"b6",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"69",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"25",x"25",x"45",x"49",x"92",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"20",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"20",x"49",x"24",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"b2",x"92",x"92",x"92",x"b2",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"92",x"b6",x"db",x"ff",x"db",x"92",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"d6",x"ff",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"49"),
     (x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"92",x"48",x"44",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"b6",x"49",x"24",x"48",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"b2",x"6d",x"69",x"49",x"49",x"49",x"49",x"69",x"92",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b2",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"20",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"45",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"45",x"24",x"24",x"49",x"45",x"49",x"25",x"24",x"49",x"92",x"49",x"49",x"25",x"25",x"25",x"b6",x"49",x"25",x"49",x"49",x"45",x"45",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"69",x"6d",x"b2",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"45",x"45",x"25",x"49",x"b6",x"24",x"25",x"45",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"20",x"24",x"00",x"20",x"20",x"20",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"45",x"92",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"92",x"69",x"49",x"6d",x"92",x"b6",x"db",x"d7",x"49",x"25",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"8e",x"ff",x"8d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b6",x"ff",x"db",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"db",x"ff",x"ff",x"db",x"92",x"49",x"6d",x"6d",x"49",x"6d"),
     (x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"92",x"6d",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"25",x"24",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"49",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"d7",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"6e",x"6d",x"49",x"49",x"49",x"25",x"24",x"92",x"49",x"49",x"49",x"49",x"25",x"49",x"6e",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"b6",x"db",x"69",x"6d",x"49",x"6d",x"49",x"6d",x"db",x"b6",x"b2",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"69",x"db",x"92",x"6d",x"6d",x"92",x"6e",x"49",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"25",x"49",x"24",x"25",x"92",x"25",x"24",x"24",x"24",x"25",x"49",x"b2",x"24",x"25",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"00",x"24",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"25",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"b2",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"69"),
     (x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"b2",x"24",x"44",x"49",x"44",x"24",x"49",x"49",x"45",x"24",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"69",x"92",x"92",x"6d",x"69",x"49",x"49",x"6d",x"b2",x"ff",x"b2",x"49",x"49",x"49",x"49",x"45",x"45",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"b2",x"92",x"92",x"b6",x"b6",x"92",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"25",x"00",x"00",x"00",x"20",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"00",x"00",x"00",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"25",x"24",x"24",x"6d",x"49",x"49",x"25",x"24",x"24",x"49",x"6d",x"49",x"49",x"45",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"6e",x"92",x"6e",x"92",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"49",x"92",x"8e",x"6d",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"45",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"00",x"00",x"20",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"b6",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"92",x"49",x"6d",x"6d",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"b6",x"49",x"44",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"92",x"6d",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"fb",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"8d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"6d",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"b6",x"92",x"6e",x"6d",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"25",x"24",x"24",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"6d",x"6d",x"45",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"6d",x"b6",x"49",x"6d",x"69",x"69",x"6d",x"92",x"ff",x"b6",x"92",x"db",x"b6",x"6d",x"6d",x"49",x"69",x"49",x"d6",x"db",x"b6",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b2",x"92",x"92",x"6e",x"6d",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"04",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"25",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"45",x"25",x"6e",x"d7",x"92",x"69",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"b2",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"db",x"db",x"fb",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"92",x"6d",x"8d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"69"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"6d",x"49",x"24",x"44",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"b6",x"92",x"6d",x"6d",x"92",x"db",x"db",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"49",x"25",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"6d",x"45",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"49",x"25",x"25",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"25",x"b6",x"49",x"49",x"49",x"49",x"45",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"6d",x"49",x"49",x"6d",x"db",x"b6",x"92",x"b2",x"b6",x"6d",x"49",x"69",x"49",x"49",x"b6",x"6d",x"49",x"6d",x"69",x"92",x"92",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"49",x"49",x"69",x"69",x"6d",x"db",x"b6",x"b6",x"92",x"b6",x"6d",x"49",x"49",x"49",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"49",x"49",x"6d",x"6d",x"25",x"49",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"92",x"db",x"b6",x"6d",x"49",x"69",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"92",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"6d",x"92",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"db",x"db",x"db",x"db",x"b6",x"b6",x"db",x"ff",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"db",x"ff",x"db",x"92",x"49",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"44",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"b6",x"92",x"b6",x"db",x"db",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"69",x"24",x"20",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"00",x"20",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"20",x"24",x"24",x"00",x"00",x"20",x"20",x"20",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"49",x"24",x"49",x"25",x"25",x"49",x"6d",x"25",x"49",x"49",x"25",x"49",x"92",x"49",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6e",x"92",x"6d",x"49",x"49",x"6d",x"6e",x"b6",x"92",x"49",x"49",x"49",x"49",x"92",x"8e",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"92",x"db",x"b2",x"b6",x"ff",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"db",x"b6",x"92",x"b6",x"db",x"49",x"6d",x"69",x"6d",x"69",x"b6",x"db",x"92",x"92",x"92",x"92",x"49",x"49",x"69",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6e",x"24",x"25",x"49",x"49",x"49",x"6d",x"24",x"25",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"20",x"49",x"45",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"45",x"45",x"45",x"49",x"69",x"92",x"d7",x"b6",x"92",x"6d",x"92",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b2",x"6d",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"45",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"b6",x"b6",x"b7",x"db",x"db",x"db",x"db",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"6d",x"48",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"45",x"45",x"45",x"24",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db",x"db",x"db",x"b6",x"92",x"8e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"25",x"25",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"69",x"6d",x"92",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"20",x"20",x"00",x"00",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"6e",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"24",x"24",x"b6",x"25",x"25",x"45",x"45",x"24",x"49",x"69",x"25",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"6d",x"d7",x"92",x"92",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"db",x"6d",x"6d",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"92",x"92",x"6d",x"69",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"72",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"20",x"00",x"20",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"45",x"49",x"49",x"8e",x"92",x"b6",x"b6",x"b6",x"b6",x"b6",x"b7",x"6e",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"44",x"24",x"24",x"24",x"69",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"fb",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"b6",x"92",x"92",x"d7",x"fb",x"fb",x"db",x"db",x"fb",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6e",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"92",x"49",x"6d"),
     (x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"6d",x"92",x"49",x"44",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"b6",x"92",x"6d",x"69",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"20",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"24",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"49",x"24",x"24",x"6d",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"6d",x"6d",x"49",x"6d",x"ff",x"b6",x"92",x"b6",x"b6",x"49",x"6d",x"49",x"49",x"49",x"db",x"b6",x"b2",x"db",x"db",x"49",x"49",x"6d",x"49",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"92",x"b6",x"92",x"b6",x"b6",x"92",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"24",x"49",x"49",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"45",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"20",x"20",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"8e",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"6d",x"92",x"6d",x"8e",x"b6",x"b6",x"db",x"db",x"b6",x"49",x"45",x"45",x"25",x"45",x"25",x"45",x"24",x"69",x"92",x"24",x"24",x"25",x"24",x"24",x"25",x"25",x"24",x"45",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"92",x"b6",x"db",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"6d",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"49",x"b6",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"92",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"25",x"49",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"25",x"6d",x"92",x"25",x"49",x"49",x"25",x"69",x"6d",x"49",x"25",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"6d",x"ff",x"b6",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"69",x"6d",x"69",x"6d",x"92",x"92",x"49",x"6d",x"49",x"49",x"b6",x"b6",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"25",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"6d",x"69",x"49",x"49",x"6d",x"92",x"b7",x"b6",x"6d",x"24",x"25",x"24",x"24",x"25",x"25",x"25",x"24",x"6d",x"6d",x"24",x"24",x"25",x"24",x"25",x"45",x"24",x"49",x"49",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"8d",x"fb",x"ff",x"ff",x"db",x"b2",x"91",x"8d",x"92",x"92",x"b6",x"db",x"92",x"92",x"8e",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"6d",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"92",x"92",x"49",x"24",x"44",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b7",x"92",x"69",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"69",x"8e",x"b6",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"8e",x"49",x"49",x"25",x"25",x"24",x"49",x"6d",x"24",x"25",x"25",x"6d",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"92",x"69",x"49",x"49",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"92",x"6d",x"69",x"6d",x"6d",x"69",x"db",x"d7",x"b6",x"b6",x"db",x"49",x"69",x"69",x"6d",x"6d",x"b6",x"92",x"6d",x"92",x"d7",x"49",x"6d",x"69",x"69",x"6d",x"ff",x"b6",x"b6",x"b6",x"db",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"6e",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"25",x"29",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"6d",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"25",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"69",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"6d",x"45",x"45",x"49",x"49",x"6d",x"92",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"25",x"24",x"24",x"45",x"45",x"45",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"b2",x"92",x"92",x"92",x"b6",x"db",x"b6",x"6e",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"b6",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"45",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"25",x"45",x"45",x"49",x"49",x"24",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"92",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"20",x"00",x"00",x"20",x"92",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"25",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"6d",x"92",x"92",x"92",x"b6",x"ff",x"6d",x"49",x"49",x"6d",x"6d",x"b6",x"6d",x"69",x"6d",x"6d",x"b6",x"6d",x"6d",x"92",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"6d",x"49",x"6d",x"b7",x"6d",x"49",x"49",x"8e",x"92",x"8e",x"92",x"b6",x"92",x"49",x"49",x"49",x"8e",x"d7",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"45",x"45",x"49",x"92",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"44",x"45",x"45",x"49",x"49",x"49",x"49",x"45",x"25",x"45",x"25",x"45",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"25",x"25",x"24",x"45",x"45",x"49",x"49",x"49",x"b2",x"db",x"8d",x"69",x"6d",x"69",x"6d",x"6d",x"6d",x"92",x"db",x"fb",x"db",x"ff",x"db",x"b6",x"92",x"92",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"24",x"92",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"8d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"6d",x"69",x"6d",x"92",x"db",x"db",x"92",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"6d",x"92",x"49",x"24",x"25",x"24",x"92",x"49",x"49",x"49",x"49",x"25",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"92",x"b6",x"69",x"6d",x"49",x"92",x"92",x"92",x"92",x"ff",x"6d",x"49",x"49",x"69",x"49",x"b6",x"92",x"6d",x"6d",x"b6",x"6d",x"49",x"69",x"49",x"6d",x"b6",x"92",x"92",x"b6",x"92",x"6d",x"69",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"ff",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"45",x"49",x"b6",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"25",x"69",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"20",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"45",x"25",x"25",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"b6",x"db",x"b7",x"db",x"fb",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6"),
     (x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"6d",x"92",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"92",x"b6",x"db",x"d7",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"49",x"6e",x"49",x"25",x"24",x"24",x"6d",x"49",x"25",x"25",x"25",x"24",x"6e",x"49",x"25",x"25",x"49",x"69",x"6e",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"69",x"6d",x"6d",x"db",x"b6",x"92",x"b6",x"db",x"6d",x"69",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"25",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b2",x"49",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b7",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"b6",x"b6",x"fb",x"db",x"db",x"d6",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"49",x"b6",x"49",x"24",x"24",x"25",x"24",x"24",x"45",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"d7",x"b6",x"d7",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"25",x"49",x"6d",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"6d",x"00",x"00",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"db",x"69",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"92",x"b6",x"92",x"b6",x"d6",x"6d",x"49",x"49",x"49",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"92",x"8d",x"b6",x"92",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"69",x"49",x"b6",x"b6",x"92",x"b6",x"ff",x"49",x"49",x"69",x"49",x"92",x"8d",x"49",x"49",x"49",x"6d",x"ff",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"49",x"69",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"24",x"49",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"92",x"b6",x"b2",x"6d",x"69",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"db",x"db",x"fb",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"ff"),
     (x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"d7",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"69",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"20",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"49",x"45",x"25",x"24",x"92",x"6d",x"49",x"49",x"49",x"25",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"92",x"db",x"b6",x"92",x"b6",x"92",x"49",x"49",x"6d",x"d6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"b6",x"ff",x"49",x"6d",x"6d",x"6d",x"6d",x"ff",x"b6",x"b6",x"db",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"49",x"92",x"db",x"92",x"92",x"b6",x"92",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"b6",x"45",x"49",x"49",x"49",x"92",x"49",x"24",x"25",x"25",x"49",x"6e",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"25",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"92",x"92",x"b6",x"92",x"92",x"92",x"92",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"b2",x"b6",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff"),
     (x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"49",x"69",x"49",x"49",x"49",x"69",x"49",x"69",x"b6",x"ff",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"25",x"49",x"25",x"49",x"49",x"25",x"6d",x"ff",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"20",x"6d",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"25",x"24",x"92",x"49",x"25",x"25",x"49",x"49",x"92",x"45",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"6e",x"92",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"49",x"92",x"db",x"b2",x"92",x"db",x"6d",x"69",x"69",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"6d",x"69",x"6d",x"ff",x"b6",x"92",x"b6",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"6e",x"24",x"25",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6e",x"6d",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"49",x"6d",x"8e",x"92",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"8d",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"fb",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"49",x"49",x"49",x"b6",x"ff",x"92",x"6d",x"69",x"6d",x"49",x"49",x"49",x"69",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"25",x"24",x"25",x"25",x"24",x"24",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"6e",x"49",x"6d",x"92",x"ff",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"db",x"92",x"db",x"b6",x"6d",x"69",x"69",x"6d",x"db",x"b6",x"b2",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"ff",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"92",x"b6",x"6e",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"69",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"6e",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"6d",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db",x"fb",x"b6",x"92",x"92",x"92",x"b2",x"b6",x"b6",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"6d",x"69",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"92",x"ff",x"db",x"6d",x"69",x"6d",x"69",x"49",x"49",x"6d",x"69",x"6d",x"db",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"45",x"49",x"49",x"25",x"49",x"8e",x"6d",x"49",x"49",x"49",x"92",x"db",x"b6",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"20",x"00",x"00",x"20",x"20",x"00",x"24",x"20",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"49",x"24",x"20",x"20",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"25",x"25",x"45",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"92",x"92",x"92",x"b6",x"db",x"49",x"49",x"6d",x"49",x"b6",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"69",x"6d",x"b6",x"92",x"6d",x"6d",x"b2",x"92",x"6d",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"92",x"92",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"6e",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"25",x"24",x"6d",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"25",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"69",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"25",x"49",x"49",x"49",x"b2",x"db",x"6d",x"49",x"49",x"49",x"69",x"69",x"6d",x"b6",x"db",x"b6",x"db",x"db",x"b6",x"b2",x"92",x"b6",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"8e",x"b6",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"b6",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"6d",x"db",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"b2",x"ff",x"db",x"6d",x"69",x"49",x"69",x"49",x"49",x"49",x"69",x"6d",x"fb",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"49",x"b6",x"45",x"24",x"44",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"25",x"45",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"6d",x"6d",x"b2",x"b7",x"92",x"69",x"45",x"45",x"25",x"24",x"25",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"20",x"24",x"49",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"20",x"00",x"00",x"24",x"20",x"20",x"20",x"00",x"24",x"20",x"24",x"20",x"6d",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"49",x"24",x"b6",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"6d",x"6d",x"b6",x"92",x"92",x"db",x"92",x"49",x"6d",x"69",x"6d",x"db",x"92",x"8d",x"b6",x"6d",x"69",x"69",x"6d",x"92",x"b6",x"92",x"b6",x"db",x"69",x"6d",x"6d",x"6d",x"db",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"ff",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"25",x"49",x"6d",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"45",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"92",x"49",x"24",x"24",x"25",x"45",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"49",x"49",x"24",x"45",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"92",x"b6",x"b6",x"92",x"b7",x"db",x"db",x"b6",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"92",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"49",x"69",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"b6",x"69",x"24",x"45",x"45",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"25",x"49",x"49",x"25",x"25",x"6d",x"b6",x"b2",x"b6",x"b6",x"92",x"6e",x"49",x"49",x"25",x"24",x"25",x"25",x"49",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"49",x"6d",x"25",x"25",x"25",x"49",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"6d",x"92",x"92",x"6d",x"b6",x"92",x"49",x"49",x"49",x"d6",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"92",x"8d",x"6d",x"6d",x"db",x"49",x"6d",x"6d",x"6d",x"db",x"b6",x"92",x"da",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"92",x"92",x"6d",x"6d",x"db",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"6d",x"6e",x"6d",x"49",x"25",x"49",x"6d",x"6d",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"45",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"ff",x"d7",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"db",x"db",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"69",x"b2",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"8e",x"92",x"49",x"44",x"49",x"45",x"24",x"49",x"25",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"45",x"24",x"25",x"24",x"25",x"49",x"92",x"db",x"d7",x"b2",x"6d",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"45",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"25",x"49",x"49",x"45",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"49",x"69",x"25",x"25",x"24",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"db",x"b6",x"6d",x"8e",x"92",x"49",x"49",x"92",x"b6",x"69",x"69",x"69",x"6d",x"db",x"6d",x"6d",x"b6",x"6d",x"49",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"49",x"6d",x"49",x"b6",x"b6",x"92",x"b6",x"db",x"6d",x"6d",x"69",x"69",x"b6",x"49",x"49",x"49",x"92",x"d7",x"92",x"92",x"92",x"6d",x"49",x"6d",x"b6",x"6e",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"25",x"49",x"92",x"49",x"24",x"25",x"49",x"49",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"49",x"49",x"45",x"24",x"24",x"00",x"24",x"20",x"00",x"20",x"24",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b2",x"6d",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"8e",x"6d",x"6e",x"b6",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"69",x"69",x"6d",x"49",x"69",x"92",x"fb",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"92",x"ff",x"db",x"8e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"92",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"45",x"49",x"49",x"25",x"45",x"49",x"24",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"b6",x"8e",x"49",x"45",x"24",x"25",x"49",x"45",x"45",x"45",x"25",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"49",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"25",x"24",x"24",x"92",x"49",x"45",x"24",x"25",x"92",x"49",x"49",x"49",x"25",x"92",x"49",x"45",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"b6",x"69",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"db",x"6d",x"6d",x"69",x"69",x"db",x"b6",x"b6",x"ff",x"6d",x"69",x"69",x"6d",x"b6",x"db",x"b6",x"db",x"92",x"6d",x"69",x"6d",x"92",x"6d",x"49",x"49",x"8d",x"b6",x"92",x"b6",x"db",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"25",x"25",x"45",x"6e",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"20",x"24",x"6d",x"6d",x"49",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"92",x"92",x"92",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"fb",x"d7",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"db",x"ff",x"fb",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"92",x"49",x"25",x"25",x"24",x"24",x"25",x"49",x"49",x"45",x"24",x"24",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"92",x"49",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"b6",x"6d",x"69",x"69",x"49",x"db",x"92",x"6d",x"92",x"92",x"49",x"49",x"92",x"92",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"b6",x"49",x"6d",x"49",x"b6",x"b6",x"92",x"d7",x"b6",x"49",x"69",x"49",x"92",x"6d",x"49",x"49",x"49",x"db",x"69",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"6d",x"49",x"45",x"49",x"6d",x"6d",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"db",x"db",x"d6",x"92",x"91",x"91",x"b6",x"b6",x"92",x"6d",x"69",x"6d",x"6d",x"b6",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"fb",x"6d",x"25",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"45",x"69",x"b6",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"20",x"20",x"00",x"00",x"49",x"49",x"24",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"49",x"92",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"b7",x"92",x"92",x"b6",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"69",x"db",x"b6",x"92",x"db",x"92",x"49",x"49",x"49",x"b6",x"92",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"db",x"b6",x"b6",x"db",x"6d",x"69",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"92",x"db",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"b2",x"b6",x"b6",x"92",x"6d",x"49",x"6d",x"69",x"6d",x"b2",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b6",x"49",x"25",x"49",x"49",x"49",x"49"),
     (x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"b2",x"69",x"49",x"49",x"49",x"69",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"49",x"24",x"25",x"45",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"20",x"20",x"20",x"24",x"25",x"49",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"20",x"49",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"20",x"20",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"92",x"49",x"24",x"25",x"24",x"92",x"24",x"25",x"24",x"49",x"6d",x"49",x"45",x"25",x"8e",x"49",x"49",x"49",x"49",x"b7",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"92",x"49",x"49",x"6d",x"b2",x"6d",x"6d",x"6d",x"b6",x"b6",x"92",x"db",x"6d",x"6d",x"6d",x"6d",x"db",x"b6",x"92",x"b6",x"6d",x"6d",x"6d",x"6d",x"b2",x"49",x"49",x"49",x"db",x"b6",x"92",x"b6",x"8e",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"49",x"49",x"6d",x"25",x"45",x"25",x"6e",x"25",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"92",x"b2",x"db",x"db",x"da",x"d6",x"db",x"b6",x"6d",x"49",x"49",x"69",x"49",x"6d",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"db",x"6d",x"24",x"49",x"49",x"49",x"49"),
     (x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"ff",x"db",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"d7",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"d6",x"ff",x"ff",x"6d",x"69",x"49",x"49",x"49",x"6d",x"49",x"69",x"d6",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"6d",x"92",x"b6",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"49",x"49",x"49",x"49",x"6e",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"92",x"92",x"92",x"8e",x"6d",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"db",x"92",x"b2",x"b6",x"49",x"6d",x"49",x"b6",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"b6",x"6d",x"69",x"49",x"49",x"db",x"92",x"b6",x"db",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6d",x"6e",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"69",x"92",x"92",x"6d",x"6d",x"92",x"db",x"fb",x"fb",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b2",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"d6",x"6d",x"6d",x"6d",x"49",x"49",x"69",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"25",x"25",x"49",x"44",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"92",x"6d",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"25",x"24",x"24",x"25",x"49",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"24",x"25",x"24",x"92",x"49",x"25",x"45",x"25",x"92",x"49",x"45",x"45",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"6d",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"b6",x"6d",x"6d",x"69",x"6d",x"db",x"92",x"db",x"b2",x"49",x"6d",x"69",x"b6",x"b6",x"92",x"db",x"6d",x"6d",x"6d",x"6d",x"ff",x"b6",x"b6",x"db",x"6d",x"69",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"8e",x"8e",x"6d",x"92",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"6e",x"25",x"49",x"49",x"92",x"49",x"25",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"49",x"25",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"25",x"25",x"45",x"49",x"49",x"6d",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"69",x"8e",x"b6",x"ff",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"25",x"49",x"49",x"25",x"45",x"49",x"49",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"6d",x"25",x"49",x"49",x"49"),
     (x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"69",x"6d",x"49",x"92",x"ff",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"49",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"72",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"25",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"92",x"24",x"25",x"49",x"49",x"92",x"45",x"45",x"25",x"92",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"d7",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"b6",x"b2",x"92",x"b6",x"6d",x"49",x"49",x"b6",x"6d",x"69",x"49",x"92",x"92",x"92",x"b6",x"92",x"49",x"6d",x"6d",x"db",x"8e",x"6d",x"b6",x"69",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"92",x"b6",x"6d",x"b6",x"92",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"24",x"25",x"45",x"6e",x"25",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"25",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"92",x"b6",x"db",x"92",x"6d",x"69",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"45",x"49",x"25",x"24",x"45",x"49",x"49",x"49",x"b6",x"92",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"24",x"49",x"49",x"49"),
     (x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"8d",x"6d",x"8d",x"6d",x"92",x"b6",x"ff",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"45",x"49",x"49",x"45",x"24",x"24",x"b6",x"49",x"49",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"45",x"24",x"24",x"49",x"6d",x"6d",x"24",x"20",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"49",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"92",x"69",x"6d",x"92",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"b6",x"92",x"db",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"b6",x"49",x"49",x"69",x"92",x"db",x"92",x"b6",x"6d",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"d7",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"25",x"24",x"25",x"92",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"20",x"24",x"20",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"69",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"d7",x"b6",x"6e",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"db",x"6d",x"24",x"49",x"45",x"24",x"24",x"49",x"49",x"24",x"69",x"d7",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"49",x"49",x"49",x"49"),
     (x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"fb",x"ff",x"ff",x"ff",x"b6",x"92",x"8d",x"8d",x"8d",x"91",x"b6",x"ff",x"db",x"db",x"db",x"b6",x"92",x"8d",x"6d",x"6d",x"92",x"d6",x"ff",x"db",x"db",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"69",x"6d",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"6d",x"25",x"49",x"24",x"25",x"45",x"25",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"b2",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"45",x"49",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"49",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"25",x"6d",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"b6",x"49",x"49",x"6d",x"b6",x"6d",x"92",x"b6",x"49",x"69",x"49",x"b6",x"49",x"49",x"69",x"db",x"b2",x"92",x"db",x"69",x"69",x"49",x"b6",x"b6",x"92",x"db",x"49",x"69",x"49",x"6d",x"db",x"92",x"b6",x"92",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"db",x"6d",x"49",x"92",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"92",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"6d",x"00",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"b6",x"b2",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"6d",x"49",x"45",x"49",x"49",x"49",x"24",x"45",x"49",x"92",x"b6",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"24",x"49",x"49"),
     (x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"91",x"92",x"92",x"b2",x"db",x"db",x"b6",x"db",x"b7",x"b6",x"92",x"92",x"8d",x"92",x"b6",x"db",x"db",x"b6",x"b7",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"db",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"6d",x"b6",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6e",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"49",x"49",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"92",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"db",x"92",x"92",x"b6",x"49",x"49",x"6d",x"92",x"69",x"69",x"6d",x"b6",x"6d",x"b2",x"92",x"49",x"69",x"69",x"b6",x"6d",x"6d",x"b6",x"69",x"69",x"6d",x"92",x"49",x"49",x"6d",x"db",x"8d",x"92",x"92",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"45",x"49",x"49",x"92",x"45",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"d7",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"92",x"92",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"49",x"d7",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"b6",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"49",x"49"),
     (x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"db",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"db",x"db",x"b6",x"92",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"92",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"b2",x"fb",x"db",x"b7",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6e",x"45",x"25",x"25",x"24",x"24",x"49",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"25",x"24",x"49",x"49",x"69",x"25",x"24",x"49",x"92",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"b6",x"92",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"db",x"92",x"b6",x"92",x"49",x"49",x"6d",x"92",x"69",x"6d",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"b6",x"49",x"49",x"49",x"db",x"92",x"92",x"b6",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"6d",x"6e",x"49",x"69",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"25",x"20",x"24",x"24",x"00",x"00",x"00",x"20",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"49",x"b6",x"49",x"49",x"24",x"45",x"49",x"49",x"24",x"45",x"25",x"6d",x"b2",x"24",x"49",x"44",x"45",x"24",x"24",x"24",x"24",x"45",x"92",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49"),
     (x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"db",x"ff",x"db",x"92",x"92",x"92",x"92",x"d7",x"db",x"b6",x"92",x"92",x"db",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"db",x"92",x"92",x"92",x"db",x"b2",x"8d",x"6d",x"8d",x"b2",x"db",x"db",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"69",x"6d",x"b6",x"fb",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"45",x"49",x"25",x"24",x"49",x"45",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"6d",x"45",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"49",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"db",x"6d",x"b6",x"92",x"49",x"49",x"92",x"6d",x"69",x"49",x"92",x"b6",x"92",x"db",x"49",x"49",x"49",x"b6",x"b6",x"92",x"db",x"49",x"49",x"49",x"b6",x"b6",x"92",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"db",x"6d",x"6d",x"6d",x"6d",x"49",x"b6",x"6d",x"49",x"49",x"92",x"49",x"49",x"45",x"49",x"6d",x"49",x"25",x"49",x"6e",x"25",x"24",x"24",x"6e",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"20",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"49",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"92",x"db",x"92",x"69",x"49",x"49",x"6d",x"6d",x"49",x"49",x"45",x"49",x"49",x"92",x"b7",x"b6",x"69",x"45",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"92",x"25",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"45",x"24",x"49",x"49",x"45",x"24",x"45",x"49",x"b6",x"49",x"49",x"45",x"44",x"44",x"24",x"24",x"45",x"24",x"69",x"b6",x"49",x"49",x"25",x"49",x"45",x"49",x"49",x"49",x"44",x"6d",x"b6",x"49",x"49"),
     (x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"db",x"db",x"db",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"92",x"b6",x"b7",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"6d",x"6d",x"92",x"db",x"92",x"92",x"92",x"92",x"db",x"db",x"92",x"6e",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b2",x"db",x"b6",x"92",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"8e",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"20",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"69",x"b6",x"92",x"92",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"92",x"b2",x"b6",x"49",x"49",x"6d",x"b6",x"6d",x"92",x"92",x"49",x"49",x"b6",x"69",x"49",x"49",x"b6",x"92",x"92",x"b2",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"25",x"45",x"49",x"92",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"45",x"25",x"25",x"24",x"49",x"49",x"49",x"6e",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"25",x"49",x"25",x"49",x"49",x"6e",x"b6",x"6d",x"25",x"45",x"49",x"49",x"49",x"25",x"24",x"49",x"b6",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"24",x"6d",x"92",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"45",x"b6",x"6d",x"49",x"49",x"45",x"24",x"49",x"49",x"49",x"49",x"45",x"b7",x"6d",x"49"),
     (x"6d",x"8d",x"6d",x"b2",x"db",x"db",x"b6",x"b6",x"db",x"ff",x"b6",x"b2",x"92",x"b6",x"db",x"db",x"92",x"92",x"6d",x"b6",x"d6",x"db",x"b6",x"d6",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"b6",x"92",x"8d",x"6d",x"6d",x"92",x"db",x"b6",x"92",x"92",x"92",x"69",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"69",x"49",x"49",x"49",x"45",x"25",x"49",x"49",x"d7",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"25",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"49",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"6d",x"49",x"25",x"24",x"6d",x"49",x"45",x"45",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"b2",x"92",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"92",x"49",x"69",x"92",x"49",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"49",x"92",x"b6",x"92",x"db",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"49",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"49",x"92",x"49",x"25",x"49",x"6d",x"49",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"6d",x"49",x"25",x"45",x"45",x"49",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"b2",x"92",x"92",x"49",x"25",x"49",x"25",x"25",x"25",x"49",x"6e",x"92",x"49",x"45",x"49",x"49",x"45",x"49",x"24",x"25",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"25",x"25",x"49",x"49",x"25",x"45",x"49",x"b6",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"6d",x"b6",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49"),
     (x"8d",x"8d",x"92",x"d6",x"fb",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"92",x"6d",x"72",x"b6",x"db",x"db",x"db",x"db",x"fb",x"b6",x"8e",x"6d",x"6d",x"6d",x"b6",x"db",x"d6",x"d6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"b6",x"92",x"92",x"92",x"b6",x"db",x"b6",x"6d",x"6d",x"92",x"92",x"69",x"49",x"49",x"49",x"6e",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"6d",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"92",x"49",x"45",x"25",x"b6",x"45",x"49",x"49",x"b2",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"6d",x"92",x"8e",x"49",x"69",x"b6",x"49",x"49",x"6d",x"db",x"92",x"db",x"6d",x"49",x"49",x"b2",x"b6",x"8e",x"b6",x"49",x"49",x"49",x"db",x"92",x"b6",x"92",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"92",x"8e",x"8e",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"25",x"49",x"45",x"92",x"24",x"25",x"24",x"6e",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"20",x"6d",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"45",x"45",x"49",x"49",x"6d",x"49",x"49",x"49",x"8e",x"b6",x"b6",x"b6",x"6d",x"25",x"25",x"25",x"24",x"25",x"24",x"49",x"92",x"6d",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"8e",x"6e",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"45",x"24",x"b6",x"69",x"49",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"45",x"d7",x"6d"),
     (x"8d",x"92",x"b6",x"fb",x"db",x"92",x"b6",x"b6",x"ff",x"db",x"b6",x"b6",x"db",x"ff",x"b7",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"fb",x"ff",x"ff",x"db",x"8e",x"6d",x"6d",x"6d",x"6d",x"db",x"db",x"db",x"ff",x"db",x"92",x"6d",x"49",x"49",x"92",x"b6",x"b6",x"b6",x"b6",x"db",x"b6",x"6d",x"49",x"6d",x"92",x"92",x"6d",x"69",x"69",x"92",x"db",x"b7",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"25",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6e",x"49",x"6d",x"69",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"92",x"69",x"92",x"49",x"49",x"92",x"69",x"49",x"49",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"db",x"6d",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"d7",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"25",x"24",x"6d",x"49",x"25",x"45",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"6d",x"49",x"45",x"49",x"49",x"6d",x"49",x"25",x"25",x"49",x"6d",x"b6",x"b6",x"6d",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"49",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"44",x"6d",x"b6",x"24",x"44",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6"),
     (x"92",x"92",x"db",x"db",x"b6",x"92",x"92",x"b6",x"ff",x"db",x"db",x"db",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"fb",x"92",x"6d",x"49",x"49",x"49",x"92",x"b6",x"db",x"db",x"db",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"6d",x"92",x"b7",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"25",x"25",x"24",x"45",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"20",x"49",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"b6",x"6d",x"6d",x"8d",x"49",x"69",x"b6",x"49",x"49",x"49",x"b6",x"6d",x"92",x"8e",x"49",x"49",x"92",x"49",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"8e",x"6d",x"49",x"49",x"b2",x"8e",x"b6",x"8e",x"49",x"49",x"8e",x"49",x"49",x"49",x"b6",x"69",x"6d",x"6d",x"49",x"49",x"92",x"49",x"25",x"49",x"92",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"6d",x"45",x"24",x"24",x"24",x"25",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"25",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"b6",x"49",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"92",x"b6",x"fb",x"b6",x"92",x"92",x"92",x"db",x"ff",x"db",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"b6",x"db",x"b2",x"6d",x"49",x"6d",x"69",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"25",x"49",x"24",x"45",x"24",x"24",x"69",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"6d",x"25",x"25",x"24",x"6d",x"49",x"49",x"24",x"6d",x"49",x"49",x"6d",x"6d",x"24",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"b6",x"92",x"6d",x"92",x"49",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"69",x"b6",x"8e",x"db",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"b6",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"24",x"24",x"24",x"92",x"24",x"24",x"25",x"6d",x"24",x"24",x"45",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"25",x"24",x"20",x"20",x"24",x"20",x"24",x"20",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"92",x"8e",x"6d",x"6d",x"49",x"24",x"24",x"25",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"b6",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"6e"),
     (x"b6",x"db",x"db",x"92",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db",x"db",x"92",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"92",x"d7",x"92",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"20",x"00",x"24",x"24",x"24",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"24",x"25",x"6d",x"25",x"49",x"25",x"92",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"6d",x"92",x"6d",x"49",x"49",x"92",x"92",x"92",x"b2",x"49",x"49",x"6d",x"b2",x"92",x"db",x"49",x"49",x"49",x"92",x"49",x"6d",x"92",x"69",x"92",x"69",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"49",x"24",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"49",x"6d",x"92",x"92",x"6e",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"45",x"24",x"45",x"24",x"24",x"24",x"45",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"44",x"49",x"b6",x"49",x"49",x"44",x"49",x"49",x"49",x"49",x"44",x"45",x"49"),
     (x"db",x"fb",x"b6",x"92",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"6d",x"69",x"69",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"b6",x"b2",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"20",x"00",x"49",x"24",x"00",x"00",x"24",x"24",x"20",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"8e",x"24",x"24",x"6d",x"49",x"24",x"24",x"92",x"24",x"24",x"49",x"69",x"45",x"45",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"6d",x"8e",x"6d",x"49",x"49",x"92",x"49",x"49",x"92",x"6d",x"6d",x"b6",x"49",x"49",x"8e",x"b2",x"8d",x"b6",x"49",x"49",x"8e",x"6d",x"49",x"92",x"6d",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"45",x"49",x"6d",x"45",x"25",x"25",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"6d",x"24",x"00",x"04",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"45",x"25",x"24",x"24",x"45",x"45",x"49",x"b6",x"49",x"45",x"24",x"24",x"24",x"49",x"24",x"44",x"44",x"6d",x"92",x"24",x"45",x"49",x"49",x"49",x"49",x"45",x"45",x"49"),
     (x"db",x"db",x"92",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"6e",x"df",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"b6",x"b6",x"69",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"49",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"6d",x"45",x"49",x"6d",x"49",x"92",x"49",x"45",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"92",x"6d",x"92",x"49",x"49",x"8e",x"49",x"49",x"8e",x"49",x"49",x"92",x"49",x"49",x"92",x"49",x"49",x"92",x"69",x"49",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"92",x"45",x"49",x"49",x"6d",x"45",x"25",x"92",x"45",x"24",x"49",x"6d",x"24",x"24",x"69",x"25",x"24",x"45",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"92",x"6d",x"25",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"92",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"25",x"49",x"92",x"6d",x"44",x"24",x"24",x"24",x"49",x"45",x"25",x"44",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25"),
     (x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"6e",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"db",x"92",x"49",x"45",x"24",x"45",x"49",x"69",x"49",x"49",x"69",x"b6",x"b6",x"6d",x"49",x"25",x"49",x"24",x"24",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"20",x"20",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"24",x"00",x"49",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"25",x"24",x"6d",x"45",x"24",x"6d",x"49",x"25",x"6d",x"92",x"49",x"6d",x"45",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"6d",x"6d",x"49",x"8e",x"49",x"49",x"92",x"6d",x"6d",x"8e",x"49",x"49",x"92",x"92",x"6d",x"92",x"49",x"49",x"6d",x"45",x"49",x"49",x"6d",x"45",x"6d",x"6d",x"69",x"6d",x"49",x"24",x"6d",x"45",x"24",x"24",x"69",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"45",x"6d",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"6d",x"92",x"24",x"24",x"25",x"25",x"25",x"49",x"45",x"45",x"69",x"b6",x"49",x"24",x"24",x"24",x"44",x"49",x"49",x"45",x"45",x"92",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"24"),
     (x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"69",x"db",x"db",x"b2",x"49",x"25",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"6d",x"b6",x"b2",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"45",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"00",x"24",x"20",x"20",x"00",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"6d",x"24",x"24",x"92",x"25",x"45",x"49",x"49",x"49",x"45",x"92",x"69",x"6d",x"49",x"45",x"92",x"49",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"6d",x"92",x"8e",x"92",x"49",x"49",x"92",x"6d",x"8e",x"6d",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"45",x"49",x"6d",x"24",x"25",x"6d",x"24",x"24",x"45",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"b2",x"49",x"45",x"49",x"49",x"45",x"25",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"45",x"49",x"44",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44"),
     (x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"92",x"b6",x"49",x"45",x"49",x"49",x"49",x"25",x"25",x"6d",x"db",x"92",x"49",x"25",x"25",x"24",x"24",x"25",x"6d",x"92",x"b6",x"b6",x"8e",x"49",x"24",x"49",x"49",x"25",x"25",x"24",x"45",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"49",x"49",x"25",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"20",x"20",x"24",x"00",x"49",x"24",x"00",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"8e",x"45",x"24",x"6d",x"49",x"6d",x"6d",x"25",x"69",x"49",x"45",x"45",x"6e",x"49",x"69",x"6d",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"6e",x"8e",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"45",x"6d",x"69",x"92",x"49",x"45",x"49",x"49",x"25",x"24",x"92",x"45",x"25",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"49",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"6d",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45"),
     (x"6d",x"69",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"6e",x"25",x"49",x"49",x"25",x"49",x"49",x"24",x"25",x"92",x"6d",x"25",x"25",x"49",x"49",x"25",x"24",x"25",x"92",x"92",x"49",x"25",x"25",x"25",x"24",x"24",x"49",x"92",x"b7",x"b6",x"6d",x"45",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"45",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"49",x"25",x"20",x"20",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"6d",x"45",x"24",x"45",x"6d",x"24",x"24",x"6d",x"24",x"24",x"6d",x"25",x"25",x"49",x"49",x"25",x"69",x"69",x"6d",x"6d",x"45",x"45",x"6d",x"45",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"8e",x"49",x"49",x"6d",x"45",x"49",x"6d",x"69",x"92",x"45",x"49",x"45",x"6d",x"45",x"6d",x"6d",x"69",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6d",x"48",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"92",x"25",x"24",x"25",x"45",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"92",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"20",x"24",x"69",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"49",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6e",x"25",x"24",x"49",x"45",x"45",x"69",x"6d",x"6d",x"6d",x"45",x"25",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"45",x"49",x"49",x"45",x"49",x"6d",x"49",x"92",x"45",x"45",x"49",x"6d",x"49",x"49",x"25",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"6d",x"49",x"25",x"49",x"25",x"24",x"45",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"00",x"24",x"49",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"45",x"24",x"25",x"25",x"45",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"6d",x"b6",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"92",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"6d",x"49",x"6d",x"45",x"24",x"6d",x"25",x"24",x"6d",x"69",x"6d",x"49",x"45",x"45",x"6d",x"49",x"6d",x"45",x"45",x"6d",x"69",x"6d",x"49",x"45",x"49",x"8e",x"69",x"6d",x"25",x"45",x"49",x"24",x"24",x"92",x"45",x"49",x"6d",x"49",x"69",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"25",x"45",x"49",x"44",x"49",x"49",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"92",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"45",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"20",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"45",x"49",x"24",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"25",x"6d",x"49",x"49",x"49",x"49",x"6d",x"25",x"24",x"6d",x"69",x"92",x"25",x"45",x"49",x"6d",x"69",x"6d",x"45",x"25",x"6e",x"69",x"92",x"25",x"24",x"49",x"24",x"24",x"6d",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"72",x"b6",x"49",x"25",x"25",x"49",x"24",x"24",x"44",x"24",x"49",x"92",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"45",x"49",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"49",x"49",x"69",x"6d",x"24",x"24",x"6d",x"49",x"6e",x"24",x"45",x"8e",x"49",x"6d",x"24",x"24",x"6d",x"49",x"45",x"6d",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"45",x"24",x"49",x"24",x"45",x"49",x"25",x"45",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"45",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"8e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"20",x"49",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"45",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"6d",x"49",x"6d",x"45",x"45",x"49",x"6d",x"69",x"49",x"24",x"24",x"69",x"49",x"49",x"25",x"49",x"24",x"24",x"45",x"69",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"20",x"24",x"49",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"24",x"49",x"49",x"45",x"45",x"69",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"92",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"69",x"24",x"24",x"49",x"45",x"69",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"49",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"45",x"49",x"49",x"49",x"45",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"45",x"24",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"45",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"45",x"69",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"24",x"6d",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"92",x"69",x"6d",x"49",x"49",x"49",x"69",x"b6",x"ff",x"db",x"6d",x"49",x"6d",x"6d",x"49",x"69",x"69",x"b6",x"ff",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"db",x"6d",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"b7",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"b6",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"25",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"69",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"45",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"44",x"24",x"24",x"24",x"25",x"69",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"6d",x"6d",x"69",x"6d",x"49",x"92",x"db",x"ff",x"b6",x"69",x"6d",x"6d",x"49",x"6d",x"69",x"92",x"ff",x"ff",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"69"),
     (x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"49",x"92",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"20",x"24",x"20",x"00",x"24",x"20",x"00",x"49",x"24",x"00",x"25",x"24",x"00",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"45",x"24",x"49",x"45",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"45",x"24",x"49",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"45",x"24",x"24",x"69",x"49",x"49",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"49",x"00",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"49",x"49",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"44",x"24",x"45",x"45",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"b6",x"6d",x"69",x"49",x"49",x"49",x"6d",x"db",x"db",x"ff",x"92",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"da",x"6d",x"6d",x"6d",x"6d",x"49",x"69",x"69",x"8e",x"fb",x"db",x"6d",x"49",x"69"),
     (x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"92",x"49",x"45",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"44",x"24",x"45",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"49",x"25",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"92",x"49",x"49",x"45",x"45",x"45",x"49",x"6d",x"b6",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"db",x"92",x"69",x"6d",x"69",x"6d",x"6d",x"b6",x"b7",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"92",x"69",x"6d"),
     (x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"92",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"92",x"49",x"24",x"24",x"45",x"25",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"25",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"25",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"20",x"24",x"25",x"20",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"49",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"49",x"25",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b6",x"6d",x"49",x"49",x"45",x"45",x"49",x"6d",x"8e",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"92",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"db",x"db",x"fb",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"6d",x"6d"),
     (x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"6d",x"6d",x"24",x"49",x"25",x"49",x"24",x"49",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"92",x"49",x"24",x"45",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"45",x"25",x"49",x"24",x"24",x"49",x"45",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"69",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"8e",x"b6",x"6d",x"49",x"45",x"49",x"49",x"49",x"6d",x"6d",x"d7",x"92",x"49",x"49",x"49",x"49",x"6e",x"6d",x"6d",x"92",x"d7",x"92",x"6d",x"6d",x"6d",x"b6",x"92",x"6e",x"92",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"b7",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"92",x"6d"),
     (x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"24",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"92",x"6d",x"49",x"24",x"24",x"49",x"45",x"24",x"49",x"24",x"92",x"49",x"25",x"25",x"24",x"49",x"49",x"49",x"49",x"92",x"6d",x"45",x"25",x"49",x"49",x"49",x"49",x"24",x"92",x"8e",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"45",x"24",x"45",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"6d",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"92",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"92",x"6d",x"6d",x"6d",x"6e",x"49",x"49",x"49",x"b6",x"db",x"92",x"8d",x"8d",x"b6",x"92",x"6d",x"6d",x"b6",x"db",x"b6",x"8d",x"6d",x"6d",x"b6",x"b6",x"92",x"b6",x"db",x"b6",x"8d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"b6",x"6d"),
     (x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"45",x"49",x"92",x"24",x"49",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"b6",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"44",x"6d",x"92",x"25",x"49",x"45",x"49",x"49",x"45",x"49",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"49",x"b2",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"20",x"20",x"24",x"20",x"20",x"24",x"20",x"24",x"24",x"24",x"45",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"25",x"49",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"6d",x"25",x"24",x"25",x"25",x"49",x"49",x"49",x"92",x"b2",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"b7",x"b6",x"92",x"6d",x"92",x"49",x"49",x"49",x"6d",x"b6",x"d7",x"b6",x"92",x"b6",x"92",x"49",x"49",x"6d",x"b6",x"db",x"b6",x"92",x"92",x"b6",x"92",x"92",x"6e",x"b6",x"db",x"b2",x"8d",x"6d",x"6d",x"92",x"db",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92"),
     (x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"6d",x"6d",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"6d",x"92",x"49",x"24",x"24",x"49",x"45",x"49",x"49",x"45",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"45",x"49",x"45",x"49",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"20",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"92",x"69",x"45",x"45",x"49",x"49",x"24",x"24",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"24",x"25",x"49",x"8e",x"d7",x"b6",x"b2",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"d7",x"db",x"92",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"b6",x"db",x"92",x"6d",x"6d",x"92",x"db",x"db",x"92",x"6d",x"91",x"92",x"db",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"ff",x"b6"),
     (x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"44",x"24",x"92",x"49",x"44",x"49",x"49",x"49",x"44",x"45",x"49",x"24",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"20",x"20",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"6e",x"b6",x"92",x"6d",x"49",x"24",x"25",x"25",x"25",x"92",x"db",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"db",x"db",x"b2",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"92",x"92",x"92",x"db",x"db",x"db",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db"),
     (x"92",x"6e",x"49",x"49",x"25",x"49",x"44",x"24",x"24",x"24",x"49",x"92",x"24",x"49",x"49",x"49",x"44",x"49",x"45",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"6e",x"92",x"6e",x"49",x"24",x"24",x"49",x"24",x"49",x"92",x"b7",x"b2",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"b2",x"b2",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff"),
     (x"b6",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"8e",x"49",x"44",x"49",x"45",x"49",x"49",x"49",x"45",x"44",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"45",x"25",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"69",x"8e",x"db",x"ff",x"b6",x"b6",x"db",x"b6",x"b2",x"92",x"b6",x"fb",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff"),
     (x"b2",x"45",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"48",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"25",x"24",x"24",x"49",x"b2",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"45",x"00",x"00",x"24",x"20",x"20",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"45",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"fb",x"db",x"db",x"db",x"b6",x"92",x"92",x"92",x"d7",x"db",x"92",x"91",x"6d",x"6d",x"92",x"d6",x"ff",x"ff"),
     (x"6d",x"25",x"44",x"24",x"49",x"49",x"24",x"24",x"48",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"fb",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"6d",x"69",x"49",x"49",x"49",x"8e",x"b6",x"6d",x"49",x"49",x"49",x"25",x"25",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"20",x"20",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"6e",x"6d",x"92",x"db",x"db",x"92",x"8d",x"8d",x"92",x"b6",x"ff",x"ff"),
     (x"49",x"25",x"45",x"49",x"49",x"49",x"44",x"49",x"24",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"b6",x"69",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"25",x"24",x"49",x"49",x"49",x"49",x"92",x"92",x"45",x"24",x"24",x"49",x"24",x"25",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"20",x"49",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"24",x"20",x"00",x"20",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"25",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"49",x"92",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"69",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6e",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff"),
     (x"25",x"25",x"44",x"49",x"49",x"48",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"69",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b7",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"8e",x"6d",x"92",x"b6",x"6d",x"25",x"24",x"24",x"49",x"6d",x"6d",x"92",x"92",x"25",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"25",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"69",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff"),
     (x"25",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"69",x"49",x"6d",x"db",x"db",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"b6",x"b6",x"6d",x"49",x"25",x"25",x"6d",x"92",x"b6",x"db",x"6d",x"25",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"6d",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"49",x"00",x"24",x"00",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b7",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b2",x"db",x"da",x"b6",x"92",x"b6",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"69",x"49",x"49",x"92",x"db",x"92",x"92",x"6d",x"69",x"69",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"b6",x"b7",x"db",x"6e",x"49",x"45",x"25",x"24",x"49",x"b6",x"db",x"92",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"45",x"20",x"20",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"00",x"24",x"20",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"6d",x"49",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"20",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"db",x"ff",x"b6",x"6d",x"49",x"69",x"6d",x"6d",x"db",x"ff",x"d6",x"b6",x"b6",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"69",x"49",x"6d",x"db",x"b6",x"6d",x"92",x"92",x"6d",x"6d",x"92",x"db",x"b2",x"49",x"49",x"49",x"49",x"92",x"db",x"fb",x"92",x"49",x"49",x"49",x"24",x"24",x"49",x"b7",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"20",x"20",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"45",x"24",x"49",x"49",x"25",x"24",x"25",x"6d",x"24",x"49",x"6d",x"25",x"25",x"49",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"49",x"b7",x"69",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"69",x"6d",x"92",x"ff",x"db",x"d6",x"d6",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"ff",x"ff",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"69",x"92",x"92",x"92",x"b2",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"45",x"49",x"49",x"25",x"25",x"6d",x"49",x"25",x"49",x"6d",x"24",x"25",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"b6",x"8e",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"ff",x"d7",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"db",x"db",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"b6",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"92",x"b6",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"45",x"49",x"b6",x"b7",x"69",x"25",x"25",x"49",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"45",x"24",x"49",x"24",x"6d",x"49",x"25",x"49",x"6d",x"49",x"49",x"49",x"6d",x"45",x"49",x"6d",x"49",x"24",x"49",x"49",x"25",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"fb",x"ff",x"db",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"92",x"d7",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"6e",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"20",x"20",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"25",x"00",x"00",x"00",x"20",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"20",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"69",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"db",x"b6",x"b6",x"6d",x"6d",x"92",x"d6",x"db",x"6d",x"49",x"49",x"49",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"24",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"ff",x"ff",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"69",x"69",x"49",x"49",x"49",x"6d",x"6d",x"db",x"db",x"b6",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6e",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"6d",x"45",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"20",x"25",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"69",x"6d",x"25",x"49",x"49",x"25",x"45",x"49",x"45",x"49",x"b6",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"6d",x"6d",x"49",x"69",x"6d",x"6d",x"b6",x"db",x"b6",x"92",x"92",x"db",x"b6",x"d6",x"fb",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"45",x"45",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"25",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"49",x"24",x"24",x"24",x"49",x"25",x"25",x"6d",x"db",x"49",x"49",x"49",x"6d",x"49",x"49",x"69",x"92",x"ff",x"ff",x"ff"),
     (x"6d",x"49",x"49",x"49",x"69",x"b6",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"b6",x"92",x"6e",x"92",x"db",x"db",x"fb",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff"),
     (x"6d",x"49",x"6d",x"69",x"6d",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"45",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"6d",x"45",x"49",x"49",x"6d",x"49",x"69",x"6e",x"69",x"6d",x"49",x"92",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"44",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"49",x"25",x"45",x"49",x"24",x"24",x"45",x"24",x"92",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"49",x"49",x"25",x"24",x"24",x"25",x"45",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff"),
     (x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"45",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6e",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"20",x"20",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"92",x"49",x"24",x"49",x"24",x"24",x"49",x"25",x"6d",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"25",x"49",x"92",x"24",x"49",x"49",x"24",x"24",x"24",x"45",x"25",x"6d",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff"),
     (x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"24",x"20",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"49",x"24",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"25",x"25",x"45",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"20",x"00",x"24",x"00",x"24",x"6e",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"d7",x"49",x"45",x"45",x"49",x"25",x"45",x"49",x"49",x"b6",x"49",x"25",x"49",x"45",x"49",x"24",x"49",x"25",x"92",x"49",x"49",x"49",x"24",x"24",x"24",x"45",x"25",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff"),
     (x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"d7",x"92",x"8d",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"92",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"20",x"20",x"20",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"45",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"6e",x"49",x"6e",x"92",x"49",x"49",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"45",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"45",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"24",x"00",x"00",x"25",x"6d",x"24",x"20",x"24",x"20",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"49",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"25",x"24",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"49",x"24",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"6d",x"25",x"49",x"49",x"24",x"24",x"25",x"45",x"25",x"b2",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff"),
     (x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"b6",x"92",x"92",x"6d",x"92",x"d6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"45",x"24",x"24",x"24",x"24",x"24",x"6e",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6e",x"6d",x"49",x"92",x"49",x"92",x"6d",x"6e",x"92",x"6d",x"8d",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"25",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"24",x"20",x"24",x"00",x"20",x"49",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"6d",x"45",x"24",x"45",x"24",x"24",x"49",x"b2",x"49",x"44",x"24",x"24",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"45",x"25",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"29",x"25",x"49",x"49",x"24",x"24",x"45",x"25",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db"),
     (x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6e",x"49",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"20",x"00",x"24",x"24",x"24",x"69",x"24",x"00",x"24",x"20",x"00",x"24",x"69",x"24",x"00",x"00",x"20",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"49",x"92",x"92",x"49",x"8e",x"92",x"92",x"92",x"49",x"92",x"49",x"49",x"92",x"6d",x"92",x"49",x"6d",x"49",x"49",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"45",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"20",x"45",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"45",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"6e",x"6d",x"49",x"49",x"24",x"24",x"24",x"6d",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"45",x"49",x"6e",x"d7",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"25",x"49",x"25",x"25",x"25",x"25",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"6d",x"92",x"b6",x"ff",x"db",x"db",x"b6",x"92",x"b2",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"45",x"6d",x"24",x"45",x"49",x"24",x"24",x"24",x"25",x"25",x"92",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"45",x"b2",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"49",x"25",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"20",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"49",x"49",x"25",x"49",x"92",x"49",x"6d",x"69",x"6d",x"49",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"92",x"6d",x"92",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"49",x"24",x"24",x"49",x"b6",x"8e",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"25",x"49",x"25",x"25",x"24",x"24",x"92",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"6d"),
     (x"6d",x"92",x"db",x"ff",x"b7",x"db",x"b6",x"b6",x"b6",x"db",x"fb",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"44",x"45",x"24",x"49",x"6d",x"24",x"45",x"49",x"24",x"24",x"25",x"25",x"49",x"8e",x"24",x"24",x"25",x"45",x"25",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"69",x"24",x"24",x"24",x"24",x"24",x"8e",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"00",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"6d",x"49",x"92",x"92",x"49",x"49",x"92",x"92",x"92",x"6d",x"92",x"49",x"92",x"92",x"49",x"92",x"6d",x"92",x"92",x"6d",x"49",x"92",x"49",x"49",x"49",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"6d",x"49",x"24",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"45",x"49",x"45",x"25",x"25",x"25",x"8e",x"69",x"25",x"24",x"49",x"24",x"45",x"49",x"49",x"49"),
     (x"6d",x"b6",x"ff",x"db",x"b6",x"db",x"b6",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"6d",x"49",x"25",x"25",x"49",x"25",x"24",x"49",x"25",x"92",x"49",x"25",x"25",x"25",x"49",x"45",x"24",x"6d",x"b6",x"45",x"24",x"24",x"24",x"25",x"45",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"45",x"24",x"24",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"92",x"6d",x"8e",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"49",x"49",x"6d",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"6d",x"b6",x"8d",x"69",x"6d",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"69",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"25",x"6d",x"92",x"25",x"24",x"49",x"24",x"25",x"45",x"49",x"24"),
     (x"92",x"b6",x"db",x"96",x"92",x"db",x"db",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"45",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"6d",x"25",x"24",x"45",x"49",x"25",x"49",x"49",x"49",x"b6",x"49",x"49",x"45",x"25",x"49",x"49",x"49",x"b6",x"92",x"45",x"24",x"49",x"49",x"45",x"6d",x"b6",x"49",x"24",x"24",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"45",x"49",x"69",x"6d",x"49",x"8d",x"6d",x"92",x"92",x"8d",x"49",x"6d",x"92",x"92",x"92",x"69",x"92",x"6d",x"92",x"6e",x"69",x"49",x"49",x"49",x"6d",x"24",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"45",x"92",x"b6",x"8e",x"6d",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"92",x"49",x"24",x"45",x"24",x"24",x"25",x"49",x"24"),
     (x"92",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"92",x"24",x"24",x"49",x"45",x"24",x"49",x"49",x"6d",x"92",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"db",x"6d",x"45",x"24",x"49",x"49",x"49",x"b6",x"69",x"24",x"24",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"6d",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"8e",x"b2",x"92",x"49",x"b2",x"92",x"92",x"6d",x"6d",x"8e",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"92",x"6d",x"49",x"25",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"6d",x"6e",x"92",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"44"),
     (x"b6",x"db",x"92",x"6d",x"6d",x"b6",x"db",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"45",x"49",x"49",x"92",x"92",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"24",x"25",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"24",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"8e",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"24",x"45",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"24",x"6d",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"6d",x"49",x"24",x"24",x"24",x"6d",x"d6",x"92",x"69",x"69",x"6d",x"6d",x"6e",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"6d",x"44",x"44",x"24",x"24",x"24",x"49",x"49"),
     (x"db",x"b6",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"24",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"92",x"49",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"8e",x"92",x"69",x"49",x"92",x"92",x"49",x"92",x"92",x"92",x"92",x"6d",x"8d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"45",x"49",x"24",x"24",x"24",x"49",x"45",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"45",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"44",x"44",x"44",x"24",x"24",x"24",x"49"),
     (x"db",x"92",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"6e",x"49",x"49",x"25",x"49",x"45",x"24",x"24",x"45",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"25",x"49",x"6d",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"8d",x"b2",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"45",x"24",x"25",x"45",x"24",x"49",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"db",x"92",x"6d",x"6d",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"45",x"24",x"24",x"24",x"49"),
     (x"b7",x"6d",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"6d",x"49",x"49",x"25",x"49",x"25",x"24",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"24",x"24",x"49",x"92",x"b6",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"25",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"69",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6e",x"49",x"92",x"92",x"8d",x"92",x"49",x"92",x"6d",x"92",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"db",x"db",x"92",x"6d",x"49",x"49",x"6d",x"db",x"92",x"69",x"49",x"6d",x"69",x"92",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"24",x"24",x"24",x"49"),
     (x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"6e",x"b6",x"49",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"00",x"20",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"45",x"69",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"69",x"69",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"6d",x"24",x"6d",x"49",x"45",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"69",x"24",x"00",x"00",x"24",x"00",x"20",x"6d",x"24",x"20",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"db",x"92",x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"69",x"69",x"6d",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"44",x"24",x"45",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"92",x"25",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"6d",x"49",x"6d",x"b6",x"6d",x"25",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"24",x"00",x"49",x"24",x"00",x"20",x"00",x"00",x"24",x"69",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"8e",x"6d",x"6d",x"6d",x"92",x"69",x"92",x"49",x"92",x"6d",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"69",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"20",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"20",x"20",x"00",x"69",x"49",x"20",x"24",x"24",x"24",x"20",x"45",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"db",x"b2",x"49",x"49",x"49",x"49",x"6d",x"d6",x"b6",x"6d",x"69",x"6d",x"6e",x"b7",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"44",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"8d",x"db",x"6d",x"49",x"49",x"6d",x"92",x"b7",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"00",x"24",x"24",x"6d",x"00",x"00",x"20",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"49",x"92",x"6d",x"6d",x"6e",x"6d",x"92",x"69",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"69",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"92",x"b2",x"49",x"25",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"6d",x"92",x"b7",x"db",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"20",x"24",x"24",x"24",x"25",x"6d",x"24",x"00",x"00",x"24",x"24",x"6d",x"24",x"00",x"00",x"20",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"49",x"92",x"49",x"49",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"45",x"69",x"25",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"25",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"20",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"00",x"20",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"92",x"49",x"24",x"49",x"49",x"49",x"69",x"b6",x"db",x"92",x"92",x"6e",x"92",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"25",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"45",x"49",x"6d",x"b2",x"db",x"92",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"20",x"20",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"45",x"24",x"49",x"24",x"6d",x"25",x"49",x"49",x"49",x"45",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"25",x"24",x"45",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"45",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"45",x"6d",x"49",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"25",x"6d",x"45",x"6d",x"49",x"6e",x"6d",x"6d",x"49",x"6d",x"25",x"49",x"49",x"49",x"45",x"6d",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"25",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"92",x"fb",x"d7",x"b6",x"92",x"92",x"92",x"b6",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49"),
     (x"25",x"49",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b2",x"49",x"49",x"49",x"49",x"6d",x"d7",x"8e",x"49",x"24",x"45",x"6d",x"b6",x"b6",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"45",x"6e",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"45",x"49",x"25",x"24",x"25",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"49",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"45",x"45",x"6d",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"45",x"49",x"49",x"6d",x"49",x"6e",x"49",x"6d",x"49",x"49",x"45",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"25",x"49",x"24",x"6d",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"b6",x"fb",x"db",x"92",x"92",x"6d",x"6d",x"db",x"b6",x"69",x"69",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49"),
     (x"25",x"49",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"69",x"49",x"49",x"6d",x"b2",x"b6",x"49",x"49",x"24",x"24",x"49",x"b6",x"6d",x"24",x"25",x"25",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"69",x"6e",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"00",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"20",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"25",x"24",x"49",x"49",x"49",x"24",x"49",x"45",x"6d",x"25",x"49",x"49",x"92",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"25",x"49",x"25",x"6d",x"49",x"49",x"49",x"25",x"6d",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"69",x"45",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"92",x"25",x"6d",x"25",x"49",x"24",x"49",x"24",x"25",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"92",x"49",x"49",x"92",x"db",x"6d",x"69",x"69",x"69",x"49",x"69",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d"),
     (x"25",x"24",x"24",x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"d7",x"b2",x"6d",x"49",x"6d",x"92",x"d7",x"6d",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"25",x"6d",x"25",x"49",x"49",x"6d",x"6d",x"6d",x"45",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"69",x"45",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"45",x"49",x"24",x"45",x"25",x"6d",x"25",x"45",x"49",x"49",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"8e",x"6e",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"24",x"49",x"49",x"25",x"6d",x"49",x"69",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"24",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"45",x"49",x"49",x"49",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"b6",x"fb",x"b6",x"49",x"49",x"49",x"6d"),
     (x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"92",x"92",x"6d",x"92",x"db",x"b2",x"49",x"49",x"49",x"24",x"24",x"25",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"25",x"6d",x"49",x"6d",x"45",x"6d",x"49",x"49",x"49",x"8e",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"69",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"45",x"49",x"69",x"49",x"6d",x"49",x"49",x"49",x"69",x"49",x"6e",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"25",x"49",x"49",x"6d",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"6d",x"49",x"49",x"49",x"92",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"b6",x"fb",x"db",x"6d",x"6d",x"6d",x"6d"),
     (x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"8e",x"b6",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"6d",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"69",x"49",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"25",x"6d",x"24",x"49",x"24",x"25",x"45",x"24",x"49",x"24",x"25",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"45",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"45",x"25",x"49",x"24",x"49",x"25",x"49",x"24",x"25",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"fb",x"6d",x"6d",x"6d",x"6d"),
     (x"24",x"24",x"24",x"24",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"8e",x"49",x"6d",x"b6",x"d7",x"ff",x"92",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"45",x"24",x"49",x"24",x"6d",x"49",x"6d",x"25",x"49",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"b6",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"69",x"49",x"8e",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"25",x"49",x"49",x"45",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"20",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"45",x"25",x"49",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"8e",x"6d",x"69",x"92",x"49",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"45",x"6d",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"69",x"92",x"44",x"24",x"24",x"24",x"25",x"6d",x"b6",x"45",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"25",x"45",x"49",x"25",x"49",x"6e",x"92",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"92",x"6d",x"6d",x"6d",x"b2",x"db",x"ff",x"b2",x"6d",x"6d",x"6d"),
     (x"24",x"24",x"25",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"49",x"6d",x"25",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"69",x"49",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"25",x"45",x"24",x"24",x"24",x"92",x"6d",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"8e",x"45",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"8e",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"8d",x"6d",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"44",x"45",x"24",x"49",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"8d",x"8d",x"6d",x"92",x"db",x"ff",x"db",x"6d",x"6d",x"6d"),
     (x"24",x"24",x"25",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6e",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"69",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"04",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"6e",x"24",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"92",x"49",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"8e",x"45",x"49",x"45",x"45",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"45",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"69",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"25",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"45",x"49",x"24",x"49",x"25",x"24",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"b2",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"45",x"49",x"6d",x"25",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"25",x"92",x"92",x"44",x"45",x"24",x"49",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"b6",x"db",x"b2",x"92",x"92",x"b6",x"db",x"fb",x"ff",x"91",x"6d",x"6d"),
     (x"24",x"49",x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"45",x"45",x"6d",x"b7",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"45",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"6d",x"49",x"92",x"49",x"6e",x"49",x"92",x"49",x"6e",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"b6",x"8e",x"92",x"6d",x"6d",x"6d",x"69",x"25",x"6d",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"49",x"49",x"25",x"6d",x"25",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"92",x"92",x"6d",x"69",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"8e",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6e",x"49",x"49",x"25",x"49",x"45",x"49",x"24",x"25",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"00",x"20",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"24",x"24",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"25",x"8e",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"45",x"6e",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"fb",x"db",x"b6",x"92",x"b6",x"db",x"db",x"ff",x"92",x"8e",x"6d"),
     (x"24",x"49",x"24",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"24",x"25",x"49",x"92",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"45",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"00",x"00",x"24",x"6d",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"6d",x"49",x"49",x"45",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"8e",x"6d",x"92",x"49",x"8e",x"49",x"92",x"8e",x"49",x"69",x"6d",x"6d",x"45",x"69",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"6d",x"8e",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"6e",x"6d",x"6d",x"6e",x"49",x"49",x"49",x"6d",x"49",x"69",x"45",x"49",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"20",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"6e",x"92",x"49",x"24",x"24",x"24",x"45",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"25",x"25",x"45",x"24",x"24",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"69",x"b7",x"ff",x"db",x"b6",x"b6",x"db",x"b6",x"db",x"db",x"92",x"8e"),
     (x"24",x"49",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"25",x"25",x"6d",x"6d",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"25",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"25",x"49",x"49",x"6d",x"45",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"92",x"6d",x"92",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"b2",x"49",x"49",x"69",x"45",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"24",x"24",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"45",x"49",x"45",x"49",x"49",x"25",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"6d",x"6d",x"69",x"49",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"24",x"49",x"25",x"45",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"45",x"24",x"25",x"49",x"25",x"49",x"69",x"45",x"69",x"49",x"49",x"8d",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"92",x"6d",x"92",x"92",x"49",x"6d",x"49",x"92",x"49",x"92",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"25",x"6d",x"25",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"00",x"24",x"00",x"20",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"69",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"25",x"24",x"49",x"49",x"d7",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"25",x"24",x"45",x"24",x"24",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"db",x"db",x"92",x"92"),
     (x"24",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"b6",x"6e",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"25",x"45",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"b2",x"92",x"45",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"20",x"24",x"24",x"24",x"24",x"6d",x"20",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"6d",x"45",x"49",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"92",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"b6",x"49",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"b6",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"45",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"25",x"6d",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"49",x"25",x"49",x"6d",x"49",x"92",x"69",x"49",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"45",x"49",x"25",x"49",x"24",x"25",x"25",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"8e",x"6d",x"92",x"8e",x"6d",x"49",x"92",x"49",x"49",x"92",x"6d",x"92",x"92",x"49",x"92",x"49",x"6d",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"25",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"24",x"00",x"24",x"6d",x"24",x"24",x"20",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"25",x"49",x"49",x"92",x"b2",x"49",x"45",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"25",x"25",x"45",x"25",x"24",x"49",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"db",x"92",x"92",x"b6",x"fb",x"b2",x"92"),
     (x"25",x"49",x"24",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"92",x"92",x"8d",x"8d",x"db",x"db",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"45",x"45",x"24",x"49",x"db",x"49",x"49",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"92",x"8e",x"6d",x"92",x"49",x"92",x"92",x"6d",x"b6",x"49",x"92",x"92",x"b6",x"92",x"92",x"49",x"6d",x"49",x"6d",x"49",x"8e",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"24",x"25",x"25",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"69",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"24",x"6d",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"69",x"49",x"b2",x"69",x"49",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"25",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"6d",x"69",x"49",x"69",x"6d",x"6d",x"92",x"49",x"92",x"49",x"6d",x"6d",x"92",x"92",x"92",x"49",x"92",x"49",x"92",x"6d",x"92",x"92",x"49",x"92",x"49",x"92",x"92",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"45",x"49",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"69",x"45",x"24",x"00",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"d7",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"6e",x"24",x"24",x"24",x"49",x"45",x"45",x"24",x"49",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"fb",x"db",x"92",x"6d",x"92",x"db",x"d6",x"92"),
     (x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"25",x"45",x"25",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"45",x"24",x"25",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"45",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"25",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"92",x"49",x"92",x"49",x"92",x"92",x"69",x"6d",x"49",x"92",x"92",x"49",x"92",x"49",x"92",x"69",x"92",x"49",x"92",x"49",x"49",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"b6",x"6d",x"92",x"6d",x"b6",x"49",x"6d",x"8d",x"49",x"49",x"6e",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"6e",x"49",x"25",x"45",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"49",x"92",x"6d",x"49",x"6d",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"69",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"8e",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"b6",x"92",x"49",x"92",x"49",x"b6",x"b6",x"49",x"92",x"49",x"92",x"6d",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"25",x"49",x"49",x"49",x"25",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"8e",x"6d",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"45",x"49",x"24",x"49",x"92",x"49",x"24",x"24",x"49",x"49",x"45",x"24",x"45",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"db",x"92"),
     (x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"b2",x"92",x"92",x"db",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"25",x"92",x"24",x"24",x"49",x"24",x"45",x"49",x"b6",x"6d",x"24",x"24",x"49",x"6d",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"25",x"6d",x"49",x"25",x"49",x"6d",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"49",x"92",x"92",x"6d",x"b6",x"92",x"92",x"92",x"49",x"b6",x"b6",x"92",x"b6",x"49",x"49",x"92",x"92",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"69",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"92",x"8d",x"b2",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"49",x"49",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"92",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"45",x"45",x"49",x"24",x"49",x"6d",x"6e",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"6d",x"92",x"69",x"6d",x"6d",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"25",x"45",x"25",x"49",x"24",x"69",x"49",x"45",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"49",x"8d",x"b6",x"6d",x"92",x"49",x"92",x"92",x"92",x"92",x"49",x"b6",x"92",x"6d",x"b6",x"49",x"92",x"69",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"45",x"6d",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"24",x"25",x"6d",x"b6",x"49",x"49",x"49",x"45",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"6d",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"db",x"92",x"6d",x"49",x"69",x"6d",x"db",x"b6"),
     (x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b2",x"92",x"6e",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"49",x"24",x"45",x"6d",x"b6",x"25",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"6d",x"25",x"25",x"49",x"6d",x"49",x"49",x"69",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"6e",x"6d",x"92",x"49",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"b2",x"49",x"92",x"49",x"92",x"8e",x"6d",x"49",x"92",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"45",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"92",x"69",x"6d",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"6e",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"92",x"6d",x"69",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"45",x"49",x"49",x"69",x"49",x"6d",x"8e",x"49",x"6d",x"92",x"92",x"b6",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"69",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"b6",x"49",x"92",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"00",x"24",x"49",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"45",x"24",x"24",x"45",x"b6",x"6d",x"49",x"49",x"45",x"25",x"49",x"b6",x"6d",x"24",x"25",x"49",x"49",x"45",x"25",x"24",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"49",x"49",x"49",x"6d",x"b6",x"db"),
     (x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"69",x"49",x"92",x"db",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"49",x"25",x"49",x"49",x"b2",x"6d",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"49",x"20",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6e",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"6e",x"6d",x"92",x"92",x"49",x"6d",x"92",x"92",x"92",x"92",x"49",x"8e",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"8e",x"49",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"92",x"69",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"8d",x"6d",x"6d",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"49",x"25",x"24",x"49",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"92",x"49",x"b2",x"92",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"92",x"49",x"6d",x"49",x"92",x"49",x"69",x"49",x"6e",x"49",x"49",x"24",x"69",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"45",x"25",x"49",x"92",x"b6",x"49",x"45",x"49",x"49",x"45",x"25",x"24",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"92",x"db"),
     (x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"6d",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"b7",x"6d",x"45",x"49",x"45",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"25",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"6d",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"d6",x"6d",x"92",x"92",x"6d",x"92",x"49",x"92",x"8d",x"92",x"49",x"6d",x"92",x"b6",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"6d",x"6d",x"49",x"b6",x"6d",x"b6",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"45",x"24",x"49",x"24",x"49",x"49",x"b6",x"49",x"92",x"b6",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"69",x"6d",x"6d",x"49",x"6d",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"49",x"92",x"49",x"8e",x"92",x"92",x"49",x"b6",x"92",x"6d",x"92",x"69",x"92",x"b6",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6d",x"24",x"49",x"25",x"49",x"24",x"25",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"20",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"25",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"69",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"db"),
     (x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"69",x"25",x"69",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"b2",x"49",x"b6",x"b6",x"69",x"b6",x"92",x"6d",x"6d",x"49",x"92",x"b6",x"49",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"8e",x"8e",x"92",x"49",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"69",x"6d",x"92",x"6e",x"6d",x"6d",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"92",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"69",x"92",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"69",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"69",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"92",x"6d",x"8e",x"92",x"6d",x"49",x"92",x"b6",x"6d",x"b6",x"6d",x"92",x"92",x"49",x"92",x"b6",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"45",x"49",x"45",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"49",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"45",x"24",x"24",x"24",x"00",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"8e",x"db",x"8d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"6e",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"49",x"49",x"49",x"49",x"6d",x"db",x"8e",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"45",x"24",x"45",x"25",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"69",x"49",x"6d",x"49",x"4d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"92",x"6d",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"69",x"92",x"8e",x"49",x"92",x"8d",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"24",x"49",x"49",x"24",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"8e",x"6d",x"6d",x"69",x"6d",x"49",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"92",x"6e",x"6d",x"92",x"49",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"b2",x"b6",x"6d",x"92",x"6e",x"b6",x"6e",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"25",x"49",x"24",x"49",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"25",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"92",x"49",x"b6",x"92",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"92",x"b6",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"b6",x"69",x"49",x"69",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"92",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"92",x"49",x"24",x"49",x"49",x"49",x"6d"),
     (x"6d",x"6d",x"db",x"6d",x"69",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"b7",x"49",x"49",x"49",x"49",x"25",x"45",x"24",x"25",x"6d",x"49",x"45",x"25",x"24",x"49",x"45",x"49",x"b6",x"92",x"49",x"49",x"49",x"92",x"b7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"45",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"b2",x"49",x"92",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"b6",x"92",x"49",x"92",x"6d",x"92",x"49",x"b6",x"6d",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"92",x"69",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"49",x"45",x"49",x"49",x"69",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"25",x"25",x"24",x"24",x"49",x"49",x"24",x"45",x"45",x"24",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"8e",x"69",x"6d",x"92",x"92",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"49",x"45",x"49",x"49",x"24",x"49",x"6d",x"69",x"6d",x"49",x"49",x"6d",x"b2",x"6d",x"6d",x"92",x"92",x"6d",x"92",x"69",x"92",x"8e",x"6d",x"49",x"92",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"92",x"49",x"92",x"6d",x"92",x"49",x"6e",x"6d",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"6e",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b7",x"8e",x"6d",x"49",x"49",x"6e",x"db",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"24",x"49",x"49",x"45",x"49",x"49",x"49",x"b6",x"92",x"24",x"24",x"49",x"25",x"24",x"49"),
     (x"6d",x"92",x"db",x"6d",x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"45",x"92",x"49",x"45",x"25",x"49",x"49",x"45",x"6d",x"db",x"49",x"49",x"49",x"6d",x"b6",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"24",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"49",x"92",x"92",x"6d",x"49",x"92",x"b6",x"49",x"6d",x"b6",x"6d",x"b6",x"6d",x"49",x"b6",x"6d",x"6d",x"49",x"92",x"92",x"49",x"6e",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"25",x"25",x"49",x"45",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"6d",x"49",x"25",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"45",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"49",x"49",x"45",x"49",x"6d",x"6d",x"b2",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"45",x"6d",x"6d",x"b6",x"49",x"49",x"92",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"92",x"69",x"49",x"49",x"92",x"6d",x"49",x"45",x"49",x"24",x"69",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"6d",x"49",x"49",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"49",x"24",x"49",x"69",x"49",x"49",x"49",x"45",x"6e",x"92",x"24",x"24",x"25",x"25",x"24",x"25"),
     (x"6d",x"b6",x"db",x"6e",x"6d",x"69",x"69",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"45",x"45",x"45",x"49",x"45",x"49",x"92",x"49",x"45",x"45",x"49",x"45",x"49",x"92",x"92",x"45",x"24",x"49",x"6d",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"6d",x"49",x"8e",x"b6",x"6d",x"92",x"b6",x"6d",x"92",x"92",x"6d",x"b6",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"49",x"6d",x"49",x"49",x"25",x"6d",x"6d",x"49",x"6d",x"92",x"69",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"69",x"49",x"24",x"25",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"45",x"6d",x"69",x"8e",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"6d",x"69",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"6d",x"92",x"8e",x"49",x"92",x"6d",x"6d",x"92",x"49",x"92",x"92",x"49",x"b6",x"92",x"49",x"92",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"25",x"49",x"49",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"25",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"24",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"24"),
     (x"6d",x"db",x"db",x"8e",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"49",x"6d",x"6e",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"92",x"92",x"49",x"92",x"92",x"49",x"92",x"6d",x"92",x"49",x"92",x"92",x"6d",x"6e",x"49",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"45",x"49",x"92",x"49",x"49",x"49",x"24",x"25",x"24",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"24",x"49",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"6d",x"6d",x"92",x"49",x"92",x"92",x"6d",x"6d",x"92",x"92",x"49",x"6d",x"72",x"6d",x"6d",x"92",x"92",x"49",x"92",x"6d",x"49",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"6d",x"45",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"20",x"24",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24"),
     (x"92",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"45",x"25",x"49",x"45",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"8d",x"92",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"45",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"25",x"49",x"92",x"49",x"6d",x"49",x"6d",x"8e",x"49",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"92",x"6d",x"6d",x"49",x"92",x"6e",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"45",x"20",x"20",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"49",x"6d",x"24",x"49",x"49",x"6e",x"24",x"49",x"49",x"49",x"6e",x"45",x"69",x"45",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"49",x"49",x"6d",x"49",x"49",x"49",x"69",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"8e",x"69",x"49",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"24",x"25",x"24",x"49",x"49",x"24",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"49",x"49",x"45",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"6e",x"49",x"92",x"49",x"92",x"49",x"6d",x"92",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"6d",x"8e",x"49",x"92",x"92",x"49",x"6d",x"49",x"92",x"49",x"49",x"25",x"6d",x"49",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24"),
     (x"92",x"ff",x"db",x"8e",x"6d",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"24",x"49",x"25",x"25",x"45",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"24",x"24",x"49",x"45",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"69",x"6d",x"92",x"49",x"92",x"8e",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"24",x"24",x"25",x"6d",x"25",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"92",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"69",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"45",x"25",x"49",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"25",x"49",x"25",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"49",x"92",x"69",x"92",x"49",x"b6",x"92",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"92",x"6d",x"49",x"6d",x"6e",x"6d",x"49",x"49",x"6d",x"49",x"49",x"25",x"6d",x"49",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"6e",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"92",x"25",x"24",x"24",x"24",x"24",x"24"),
     (x"b6",x"ff",x"db",x"92",x"6d",x"92",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"45",x"45",x"44",x"24",x"49",x"49",x"b6",x"8e",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"20",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"45",x"25",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"92",x"8e",x"6d",x"49",x"6d",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"49",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"25",x"45",x"49",x"92",x"6d",x"45",x"92",x"49",x"45",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"25",x"45",x"24",x"45",x"45",x"49",x"69",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"45",x"24",x"49",x"45",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"49",x"8e",x"6d",x"69",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"25",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"24",x"00",x"00",x"25",x"49",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24"),
     (x"db",x"ff",x"db",x"b6",x"92",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"69",x"49",x"49",x"45",x"49",x"49",x"45",x"49",x"49",x"db",x"8e",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"25",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"25",x"49",x"25",x"49",x"6d",x"92",x"49",x"49",x"49",x"6e",x"92",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6e",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"45",x"24",x"49",x"24",x"25",x"45",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"69",x"49",x"92",x"49",x"92",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"24",x"92",x"24",x"24",x"92",x"49",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"6d",x"69",x"49",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"b6",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"24",x"25",x"25",x"6d",x"25",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"24",x"24",x"00",x"20",x"24",x"00",x"20",x"24",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"25",x"6e",x"db",x"6d",x"49",x"49",x"6d",x"92",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24"),
     (x"ff",x"ff",x"ff",x"b6",x"b6",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"49",x"49",x"45",x"45",x"49",x"49",x"49",x"6d",x"db",x"6e",x"69",x"49",x"49",x"b2",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"6e",x"6d",x"49",x"6d",x"49",x"6d",x"45",x"6d",x"25",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6d",x"92",x"49",x"69",x"49",x"92",x"49",x"25",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"69",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"49",x"25",x"49",x"45",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6e",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"45",x"49",x"25",x"6d",x"49",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"45",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"6d",x"24",x"20",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"25",x"49",x"db",x"b6",x"6d",x"69",x"6d",x"b2",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24"),
     (x"ff",x"db",x"db",x"db",x"d6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"49",x"92",x"b7",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"20",x"24",x"24",x"25",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"25",x"24",x"20",x"24",x"24",x"24",x"00",x"25",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"92",x"49",x"25",x"25",x"49",x"6e",x"69",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"45",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"b6",x"92",x"49",x"6d",x"24",x"6d",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"49",x"24",x"92",x"b6",x"49",x"92",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"25",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"25",x"92",x"db",x"92",x"8e",x"8e",x"92",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24"),
     (x"ff",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"25",x"49",x"25",x"45",x"49",x"49",x"49",x"db",x"92",x"49",x"6d",x"92",x"b6",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"25",x"20",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"45",x"25",x"6e",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"24",x"6d",x"45",x"92",x"6d",x"49",x"49",x"6d",x"69",x"49",x"25",x"25",x"24",x"20",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6e",x"49",x"69",x"49",x"6d",x"49",x"45",x"24",x"25",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"00",x"24",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"25",x"69",x"db",x"b6",x"b6",x"6e",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24"),
     (x"db",x"92",x"92",x"b6",x"db",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"db",x"6d",x"49",x"49",x"92",x"db",x"b6",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"45",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"25",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"25",x"25",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6e",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"69",x"49",x"6d",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"6d",x"24",x"49",x"92",x"92",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"25",x"6d",x"25",x"49",x"25",x"b6",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"49",x"6d",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"45",x"45",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6e",x"6d",x"25",x"49",x"24",x"6d",x"25",x"25",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"25",x"24",x"24",x"25",x"25",x"20",x"00",x"49",x"00",x"24",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"45",x"45",x"49",x"b6",x"db",x"b6",x"6d",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24"),
     (x"b7",x"6d",x"6d",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"25",x"25",x"6d",x"b6",x"6d",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6e",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"6d",x"49",x"25",x"25",x"25",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"25",x"49",x"6d",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"6d",x"b6",x"24",x"6e",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"45",x"24",x"25",x"24",x"49",x"6d",x"24",x"6d",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"49",x"24",x"49",x"24",x"49",x"6d",x"25",x"6d",x"49",x"45",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"6d",x"24",x"45",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"25",x"6d",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"49",x"49",x"b6",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"45",x"49",x"25",x"6d",x"b6",x"92",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"49",x"24",x"24"),
     (x"92",x"6d",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8e",x"25",x"24",x"24",x"49",x"92",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"24",x"24",x"20",x"24",x"45",x"20",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"25",x"6d",x"49",x"6d",x"49",x"49",x"69",x"6d",x"49",x"49",x"6d",x"6d",x"45",x"49",x"49",x"6d",x"25",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"24",x"92",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"92",x"49",x"6d",x"24",x"49",x"69",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"6d",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"69",x"49",x"24",x"49",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"25",x"45",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"24",x"24"),
     (x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"24",x"24",x"24",x"49",x"72",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"69",x"b6",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"00",x"20",x"24",x"20",x"20",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"45",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"69",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"25",x"6e",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"25",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"25",x"24",x"49",x"49",x"24",x"25",x"6e",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"25",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"00",x"24",x"49",x"24",x"00",x"24",x"49",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"24",x"24",x"20",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"24",x"24"),
     (x"49",x"49",x"49",x"49",x"8e",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"20",x"20",x"49",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"25",x"24",x"49",x"49",x"6e",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"49",x"6d",x"49",x"25",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"69",x"24",x"24",x"6d",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"25",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"69",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"6e",x"49",x"25",x"24",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"49",x"49",x"49",x"49",x"45"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"6e",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"6d",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"25",x"45",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"25",x"45",x"49",x"49",x"24",x"69",x"49",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"69",x"92",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"20",x"24",x"49",x"24",x"24",x"20",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"25",x"69",x"db",x"6d",x"49",x"49",x"49",x"49",x"69",x"b6",x"6d",x"49",x"49",x"49",x"49"),
     (x"49",x"25",x"24",x"49",x"6d",x"b2",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"20",x"00",x"25",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"45",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"8e",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"6d",x"49",x"24",x"25",x"49",x"45",x"49",x"b6",x"92",x"69",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49"),
     (x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"69",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"92",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"45",x"49",x"24",x"25",x"49",x"24",x"49",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"20",x"24",x"49",x"00",x"20",x"49",x"00",x"00",x"25",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"49",x"24",x"25",x"49",x"49",x"45",x"92",x"d6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49"),
     (x"24",x"24",x"24",x"24",x"6d",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"6d",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"45",x"25",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"00",x"49",x"24",x"00",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"69",x"25",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"92",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"25",x"25",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"69",x"24",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"25",x"49",x"6d",x"b2",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"45",x"6d",x"db",x"92",x"6d",x"69",x"49",x"6d",x"b6",x"db",x"69",x"49",x"49",x"49"),
     (x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b2",x"6d",x"6d",x"6d",x"b6",x"db",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"b6",x"49",x"49",x"49",x"6d",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"6d",x"20",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"49",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"25",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"69"),
     (x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"8e",x"ff",x"92",x"6d",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"25",x"25",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"49",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"92",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"24",x"69",x"49",x"24",x"24",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"45",x"49",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"24",x"00",x"20",x"00",x"49",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"45",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"92",x"db",x"ff",x"6d",x"49",x"69",x"6d"),
     (x"24",x"24",x"24",x"24",x"69",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"6d",x"92",x"db",x"ff",x"6e",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"25",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"49",x"24",x"49",x"49",x"25",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"49",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"49",x"20",x"20",x"49",x"00",x"00",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"45",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"92",x"6d",x"6d",x"69"),
     (x"24",x"24",x"24",x"24",x"69",x"69",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"6e",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"b6",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"45",x"24",x"6d",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"69",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"45",x"24",x"49",x"24",x"6d",x"24",x"6d",x"24",x"49",x"49",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"69",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"00",x"45",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"6d",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"72",x"49",x"49",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"45",x"49",x"49",x"49",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"92",x"6d",x"6d",x"69"),
     (x"24",x"24",x"24",x"24",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"6d",x"6d",x"92",x"db",x"b7",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"25",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"69",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"db",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"49",x"6d",x"92",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"69",x"49",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"20",x"20",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"45",x"45",x"49",x"49",x"49",x"49",x"b6",x"db",x"db",x"b6",x"92",x"b6",x"ff",x"b6",x"6d",x"6d",x"69"),
     (x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"44",x"b2",x"69",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"20",x"49",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"24",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"49",x"b2",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"25",x"00",x"20",x"00",x"45",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"49",x"b7",x"49",x"25",x"45",x"49",x"24",x"24",x"49",x"49",x"24",x"45",x"45",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"92",x"8e",x"92",x"db",x"db",x"6d",x"69",x"69"),
     (x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"6d",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"6d",x"25",x"24",x"45",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"25",x"49",x"45",x"6d",x"24",x"25",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"45",x"24",x"25",x"24",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"b6",x"25",x"92",x"49",x"8d",x"69",x"49",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"92",x"24",x"49",x"49",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"6d",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"8e",x"92",x"6d",x"92",x"6d",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"92",x"45",x"49",x"25",x"25",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"69",x"24",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"20",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"24",x"45",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"6d",x"92",x"b6",x"db",x"6d",x"49",x"69"),
     (x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"25",x"49",x"6e",x"6d",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"6d",x"25",x"24",x"25",x"44",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"49",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"49",x"20",x"00",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"6d",x"24",x"24",x"69",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"69",x"24",x"49",x"49",x"24",x"6d",x"24",x"6d",x"49",x"49",x"49",x"45",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"6d",x"49",x"6d",x"92",x"92",x"25",x"49",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"6d",x"25",x"49",x"24",x"25",x"49",x"24",x"92",x"49",x"69",x"6d",x"25",x"49",x"6d",x"6d",x"45",x"25",x"24",x"24",x"69",x"49",x"6d",x"24",x"6d",x"6d",x"92",x"6d",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"25",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"6d",x"24",x"69",x"24",x"49",x"69",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"25",x"49",x"49",x"49",x"6d",x"24",x"25",x"49",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"8e",x"92",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"24",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"8d",x"49",x"49"),
     (x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"b7",x"6d",x"25",x"25",x"25",x"25",x"6d",x"49",x"25",x"49",x"49",x"25",x"49",x"24",x"25",x"92",x"92",x"49",x"25",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"69",x"25",x"69",x"69",x"6d",x"49",x"6e",x"49",x"49",x"6d",x"24",x"69",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"49",x"6d",x"6d",x"45",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"8e",x"49",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"92",x"24",x"49",x"24",x"24",x"49",x"6d",x"49",x"24",x"45",x"49",x"6d",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"69",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"25",x"45",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"25",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"6d",x"24",x"24",x"69",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"25",x"25",x"49",x"92",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"6d",x"db",x"92",x"49",x"49"),
     (x"49",x"24",x"45",x"24",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"24",x"49",x"24",x"25",x"6d",x"49",x"25",x"49",x"25",x"25",x"49",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"92",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"25",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"45",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"8e",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"69",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"24",x"6d",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"69",x"6d",x"49",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"6e",x"6d",x"6d",x"24",x"69",x"24",x"24",x"25",x"49",x"25",x"49",x"69",x"49",x"6d",x"49",x"49",x"92",x"49",x"b6",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"45",x"25",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"69",x"49",x"49",x"6d",x"6d",x"45",x"6d",x"49",x"24",x"6d",x"24",x"25",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"24",x"25",x"49",x"92",x"24",x"45",x"25",x"25",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49"),
     (x"49",x"25",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"24",x"49",x"db",x"92",x"49",x"6d",x"6d",x"b6",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"69",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"25",x"45",x"49",x"45",x"92",x"45",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"20",x"20",x"25",x"00",x"24",x"00",x"24",x"00",x"45",x"20",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"45",x"24",x"25",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"92",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"6d",x"24",x"69",x"49",x"6d",x"49",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"b6",x"49",x"49",x"45",x"44",x"6d",x"b2",x"49",x"45",x"24",x"49",x"49",x"24",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"d6",x"69",x"49"),
     (x"49",x"49",x"49",x"25",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"25",x"49",x"db",x"6d",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"45",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"69",x"24",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"25",x"6d",x"45",x"49",x"92",x"69",x"49",x"49",x"92",x"25",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"6d",x"6d",x"6e",x"6d",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"49",x"45",x"6d",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"45",x"24",x"45",x"45",x"45",x"25",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"45",x"6d",x"45",x"45",x"6d",x"45",x"6d",x"25",x"25",x"49",x"25",x"69",x"24",x"25",x"6d",x"24",x"45",x"6d",x"24",x"49",x"45",x"6d",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"20",x"20",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"49",x"49",x"24",x"25",x"45",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"45",x"49",x"25",x"49",x"db",x"49",x"25",x"49",x"6d",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"49",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"45",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"69",x"6d",x"49",x"49",x"6d",x"24",x"6d",x"45",x"45",x"69",x"45",x"49",x"45",x"25",x"6d",x"25",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"69",x"45",x"6d",x"24",x"6d",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"92",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6e",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"25",x"6d",x"24",x"6d",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"44",x"6d",x"24",x"25",x"6d",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"8e",x"b6",x"49",x"44",x"24",x"49",x"49",x"25",x"25",x"25",x"6e",x"6d",x"25",x"49",x"49",x"49",x"49",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"8e",x"db",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"6d",x"24",x"24",x"6d",x"25",x"45",x"49",x"45",x"69",x"49",x"49",x"92",x"49",x"69",x"6d",x"6d",x"24",x"8e",x"24",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"45",x"49",x"25",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"45",x"49",x"49",x"69",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"45",x"6d",x"45",x"45",x"49",x"49",x"6d",x"45",x"49",x"45",x"45",x"92",x"45",x"6d",x"49",x"8e",x"49",x"45",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"24",x"25",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"92",x"b6",x"6d",x"49",x"49",x"8e",x"b6",x"6d",x"45",x"24",x"49",x"49",x"45",x"25",x"24",x"6d",x"69",x"24",x"49",x"49",x"49",x"49",x"b6",x"92",x"49"),
     (x"49",x"49",x"49",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"45",x"24",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"25",x"00",x"00",x"24",x"00",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"25",x"49",x"24",x"6d",x"45",x"45",x"6d",x"45",x"25",x"6d",x"45",x"49",x"6d",x"49",x"6d",x"6d",x"8e",x"45",x"6d",x"45",x"45",x"49",x"45",x"69",x"45",x"6d",x"49",x"6d",x"49",x"45",x"49",x"45",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"25",x"6d",x"24",x"6d",x"6d",x"45",x"6d",x"49",x"49",x"6e",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"45",x"24",x"25",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"69",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"25",x"8e",x"24",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"92",x"45",x"49",x"49",x"45",x"6d",x"45",x"45",x"49",x"45",x"8e",x"49",x"49",x"6d",x"49",x"69",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b7",x"92",x"6d",x"69",x"8e",x"b7",x"92",x"49",x"25",x"25",x"49",x"49",x"25",x"24",x"6d",x"49",x"24",x"25",x"49",x"49",x"49",x"92",x"b6",x"6d"),
     (x"49",x"49",x"49",x"69",x"db",x"92",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"29",x"49",x"6d",x"6d",x"45",x"25",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"6d",x"24",x"24",x"49",x"25",x"25",x"92",x"45",x"49",x"8e",x"6d",x"6d",x"45",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"69",x"8e",x"6d",x"6d",x"92",x"45",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"45",x"24",x"49",x"45",x"49",x"49",x"6d",x"49",x"49",x"49",x"8e",x"49",x"6d",x"6d",x"49",x"24",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"6d",x"49",x"b6",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"6d",x"49",x"24",x"45",x"49",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"45",x"6d",x"24",x"6d",x"45",x"6d",x"45",x"49",x"45",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"69",x"49",x"49",x"45",x"45",x"6d",x"24",x"24",x"8e",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"6d",x"6e",x"b6",x"b2",x"49",x"25",x"25",x"49",x"45",x"49",x"24",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"db",x"6d"),
     (x"49",x"49",x"49",x"6d",x"db",x"92",x"69",x"49",x"6d",x"92",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"45",x"25",x"49",x"49",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"69",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"8e",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"20",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"6d",x"24",x"24",x"69",x"24",x"24",x"6d",x"49",x"69",x"6d",x"49",x"92",x"45",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"45",x"6d",x"45",x"69",x"45",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"45",x"24",x"24",x"45",x"25",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"69",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"25",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"8e",x"49",x"92",x"6d",x"69",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"69",x"45",x"8e",x"6d",x"6d",x"49",x"92",x"49",x"45",x"6d",x"25",x"25",x"6d",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"45",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6e",x"92",x"6e",x"49",x"69",x"92",x"b6",x"49",x"45",x"49",x"49",x"25",x"49",x"24",x"6d",x"49",x"24",x"45",x"45",x"49",x"49",x"49",x"db",x"92"),
     (x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"69",x"6d",x"d6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"d7",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"45",x"92",x"49",x"45",x"6d",x"49",x"49",x"6d",x"49",x"8e",x"92",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"6d",x"6d",x"8e",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"45",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"69",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"6d",x"45",x"6d",x"45",x"6d",x"49",x"6e",x"6d",x"6d",x"6d",x"b2",x"49",x"49",x"69",x"49",x"6d",x"49",x"49",x"92",x"45",x"6d",x"69",x"92",x"49",x"45",x"6d",x"45",x"25",x"6d",x"24",x"24",x"6d",x"24",x"25",x"45",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"6d",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"db",x"b2"),
     (x"49",x"49",x"69",x"92",x"ff",x"b6",x"92",x"92",x"92",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"92",x"25",x"25",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"8e",x"8e",x"92",x"49",x"6d",x"49",x"49",x"45",x"45",x"49",x"45",x"69",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"25",x"24",x"24",x"45",x"49",x"92",x"6d",x"92",x"92",x"49",x"69",x"b6",x"6d",x"6d",x"b6",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"69",x"24",x"24",x"24",x"49",x"6d",x"24",x"6d",x"49",x"24",x"49",x"49",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"69",x"6d",x"49",x"6d",x"92",x"92",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"49",x"8e",x"92",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"8e",x"49",x"6d",x"49",x"45",x"6d",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"49",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"25",x"49",x"db",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"6d",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"b6",x"b6"),
     (x"49",x"49",x"69",x"92",x"ff",x"db",x"b6",x"b6",x"b6",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"45",x"49",x"24",x"8e",x"24",x"24",x"49",x"45",x"45",x"b6",x"6d",x"6e",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"b2",x"8e",x"6d",x"6e",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"69",x"49",x"49",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"8e",x"69",x"45",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"92",x"6d",x"49",x"24",x"49",x"92",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"49",x"49",x"45",x"24",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"69",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"49",x"69",x"49",x"25",x"49",x"45",x"49",x"45",x"92",x"49",x"92",x"92",x"6d",x"69",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"6e",x"6d",x"6e",x"49",x"6d",x"49",x"49",x"49",x"45",x"45",x"92",x"49",x"49",x"49",x"24",x"6d",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"25",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"45",x"49",x"24",x"6d",x"49",x"24",x"25",x"49",x"49",x"49",x"25",x"92",x"db"),
     (x"49",x"49",x"49",x"b6",x"ff",x"db",x"b7",x"db",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"b7",x"45",x"24",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"92",x"24",x"24",x"49",x"45",x"45",x"92",x"69",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"92",x"49",x"49",x"6d",x"49",x"b6",x"6e",x"6d",x"6d",x"49",x"49",x"6d",x"45",x"6d",x"25",x"49",x"6d",x"24",x"6d",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"6e",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"6d",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"d7",x"49",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"45",x"25",x"49",x"49",x"24",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"b6",x"6d",x"6d",x"49",x"92",x"45",x"49",x"6d",x"24",x"24",x"8e",x"45",x"49",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"49",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"25",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"45",x"49",x"25",x"8e",x"49",x"24",x"25",x"49",x"49",x"49",x"45",x"6d",x"ff"),
     (x"49",x"49",x"49",x"b6",x"db",x"b6",x"92",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"92",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"25",x"6e",x"49",x"6d",x"49",x"45",x"8e",x"49",x"49",x"92",x"49",x"92",x"92",x"b6",x"49",x"49",x"6d",x"49",x"92",x"49",x"92",x"8e",x"b6",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"6d",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"8e",x"69",x"49",x"49",x"69",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"b6",x"49",x"b6",x"6d",x"49",x"8e",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"8e",x"6d",x"92",x"b6",x"49",x"8e",x"49",x"49",x"6d",x"49",x"92",x"92",x"6d",x"49",x"b6",x"49",x"49",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"92",x"49",x"25",x"6d",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"49",x"24",x"45",x"49",x"49",x"45",x"25",x"49",x"ff"),
     (x"49",x"49",x"49",x"db",x"db",x"92",x"6d",x"92",x"b7",x"fb",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"6d",x"49",x"49",x"49",x"24",x"8e",x"49",x"49",x"6d",x"49",x"6d",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"b6",x"6d",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"8e",x"6d",x"49",x"92",x"49",x"49",x"45",x"8e",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"25",x"24",x"6d",x"25",x"6e",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"69",x"6d",x"49",x"49",x"24",x"24",x"25",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"49",x"24",x"6d",x"24",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"b2",x"69",x"92",x"92",x"92",x"49",x"92",x"49",x"49",x"92",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"24",x"6d",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"45",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"49",x"49",x"49",x"45",x"25",x"49",x"db"),
     (x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"69",x"b6",x"db",x"49",x"25",x"49",x"49",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"20",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"92",x"25",x"25",x"6d",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"6d",x"92",x"49",x"92",x"49",x"49",x"92",x"49",x"92",x"b2",x"8e",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"45",x"6d",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"69",x"6d",x"25",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"45",x"49",x"6d",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"6e",x"24",x"25",x"24",x"25",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"6d",x"6e",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"45",x"25",x"49",x"69",x"25",x"6d",x"92",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"45",x"49",x"45",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"92",x"49",x"8e",x"49",x"6d",x"b2",x"db",x"49",x"69",x"6d",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"b7"),
     (x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"6d",x"db",x"db",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"6d",x"24",x"24",x"49",x"45",x"45",x"6e",x"6d",x"92",x"49",x"49",x"92",x"49",x"49",x"b2",x"92",x"6d",x"49",x"92",x"49",x"6d",x"6d",x"8d",x"92",x"b6",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"8e",x"49",x"49",x"49",x"6d",x"49",x"69",x"49",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"45",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"92",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"25",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"45",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"6d",x"24",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"49",x"92",x"92",x"6d",x"b6",x"49",x"49",x"6d",x"49",x"b6",x"92",x"6d",x"49",x"b6",x"49",x"49",x"92",x"49",x"92",x"6d",x"b6",x"49",x"49",x"6d",x"25",x"49",x"92",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"b2"),
     (x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"6d",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"6e",x"b7",x"b6",x"25",x"25",x"49",x"24",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"25",x"49",x"b6",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"6d",x"25",x"24",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"b6",x"6d",x"92",x"49",x"92",x"49",x"49",x"b2",x"49",x"92",x"6d",x"b6",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"69",x"25",x"45",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6d",x"25",x"6d",x"45",x"92",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"b6",x"49",x"b6",x"92",x"6d",x"49",x"92",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"b6",x"49",x"49",x"6d",x"24",x"24",x"6d",x"25",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"04",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92"),
     (x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"6d",x"92",x"b6",x"92",x"25",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"25",x"49",x"6e",x"b6",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"6d",x"45",x"25",x"49",x"45",x"8e",x"49",x"49",x"92",x"49",x"6d",x"49",x"69",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"49",x"92",x"49",x"92",x"6d",x"b6",x"49",x"6d",x"49",x"92",x"8d",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"45",x"6d",x"24",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"25",x"6d",x"6d",x"6d",x"6e",x"49",x"92",x"49",x"92",x"6d",x"92",x"6d",x"92",x"49",x"92",x"49",x"92",x"92",x"b6",x"49",x"6d",x"49",x"49",x"b6",x"6d",x"6d",x"49",x"8d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"24",x"25",x"6d",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"25",x"24",x"24",x"25",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"b2",x"69",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"92"),
     (x"49",x"49",x"6e",x"d7",x"49",x"49",x"25",x"29",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"49",x"92",x"6e",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"92",x"45",x"49",x"6d",x"49",x"49",x"6d",x"49",x"b6",x"49",x"49",x"92",x"49",x"92",x"69",x"b6",x"49",x"49",x"b2",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"8e",x"6d",x"45",x"49",x"25",x"49",x"49",x"25",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"25",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"45",x"49",x"49",x"6d",x"92",x"49",x"92",x"49",x"92",x"49",x"92",x"92",x"b6",x"69",x"6d",x"49",x"49",x"db",x"b6",x"6d",x"49",x"92",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6e",x"24",x"24",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"00",x"20",x"00",x"00",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"45",x"49",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"db",x"92",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"8e"),
     (x"49",x"49",x"92",x"b6",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"24",x"49",x"6d",x"6d",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"92",x"6d",x"45",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"6d",x"49",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"49",x"92",x"49",x"6d",x"92",x"b6",x"49",x"49",x"92",x"49",x"92",x"b6",x"49",x"49",x"8e",x"49",x"92",x"b2",x"49",x"49",x"49",x"6d",x"69",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"6e",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"25",x"45",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"45",x"24",x"24",x"25",x"49",x"25",x"49",x"25",x"6d",x"6d",x"92",x"49",x"49",x"49",x"92",x"6d",x"6d",x"b6",x"49",x"6d",x"69",x"69",x"b6",x"db",x"49",x"49",x"6d",x"49",x"92",x"8d",x"92",x"49",x"49",x"6d",x"49",x"92",x"6d",x"92",x"49",x"49",x"92",x"49",x"49",x"92",x"49",x"6d",x"24",x"24",x"6d",x"24",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"6d"),
     (x"49",x"49",x"b2",x"92",x"49",x"25",x"49",x"49",x"25",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"25",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"20",x"24",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"6d",x"24",x"25",x"49",x"6e",x"49",x"6d",x"49",x"6e",x"49",x"49",x"92",x"92",x"d7",x"49",x"49",x"92",x"49",x"92",x"92",x"db",x"49",x"6d",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"92",x"92",x"6d",x"92",x"49",x"92",x"49",x"6d",x"6d",x"45",x"49",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"45",x"24",x"24",x"92",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"25",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"92",x"24",x"92",x"49",x"24",x"6d",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"45",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"b6",x"b6",x"49",x"49",x"8d",x"49",x"b6",x"92",x"92",x"49",x"92",x"49",x"49",x"b6",x"b6",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"92",x"24",x"24",x"6d",x"25",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"6d",x"44",x"25",x"25",x"24",x"49",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"92",x"db",x"6d",x"49",x"69",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"24",x"45",x"25",x"6d"),
     (x"49",x"49",x"b6",x"6d",x"49",x"25",x"49",x"49",x"24",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"b6",x"6d",x"6d",x"49",x"8e",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"92",x"49",x"92",x"6d",x"b6",x"49",x"6d",x"6d",x"92",x"49",x"92",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"25",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"24",x"25",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"92",x"92",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"6d",x"49",x"24",x"49",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6e",x"92",x"92",x"49",x"8e",x"49",x"b6",x"92",x"8e",x"49",x"92",x"49",x"92",x"92",x"b6",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"25",x"45",x"92",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"25",x"49",x"45",x"8e",x"db",x"92",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"6d"),
     (x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"b7",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"69",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"49",x"6d",x"45",x"45",x"92",x"49",x"6d",x"49",x"92",x"49",x"49",x"92",x"92",x"b6",x"49",x"49",x"92",x"49",x"92",x"92",x"92",x"49",x"92",x"69",x"92",x"49",x"92",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"45",x"49",x"25",x"69",x"69",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"25",x"45",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"6d",x"49",x"92",x"6d",x"b6",x"49",x"92",x"49",x"92",x"92",x"b6",x"49",x"6d",x"49",x"49",x"b2",x"b6",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"b6",x"49",x"49",x"45",x"45",x"6d",x"24",x"24",x"6d",x"25",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"00",x"20",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"25",x"25",x"49",x"6d",x"25",x"25",x"25",x"24",x"25",x"45",x"45",x"6d",x"b6",x"b6",x"92",x"8e",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"6d"),
     (x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"45",x"20",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"6e",x"6e",x"92",x"49",x"49",x"92",x"49",x"8e",x"49",x"92",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"92",x"49",x"92",x"6d",x"92",x"49",x"b6",x"92",x"92",x"49",x"6d",x"49",x"6d",x"8e",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"69",x"b6",x"6d",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"45",x"24",x"25",x"25",x"25",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"b6",x"49",x"92",x"49",x"92",x"92",x"92",x"69",x"8d",x"49",x"6d",x"b6",x"db",x"49",x"49",x"92",x"49",x"6d",x"49",x"b6",x"49",x"49",x"b6",x"6d",x"69",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"92",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"25",x"49",x"6d",x"92",x"49",x"45",x"45",x"24",x"25",x"25",x"45",x"49",x"92",x"b6",x"92",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d"),
     (x"49",x"8d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"49",x"25",x"44",x"49",x"24",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"6d",x"44",x"25",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"49",x"92",x"92",x"b2",x"49",x"49",x"6d",x"6d",x"92",x"92",x"6d",x"69",x"b6",x"92",x"92",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"49",x"6d",x"69",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"6d",x"92",x"45",x"25",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"92",x"b6",x"49",x"6d",x"49",x"6d",x"b6",x"d6",x"49",x"6d",x"6d",x"49",x"92",x"b6",x"6d",x"49",x"92",x"6d",x"92",x"49",x"49",x"6d",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"6d",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"6d",x"92",x"49",x"45",x"45",x"24",x"24",x"25",x"25",x"49",x"92",x"92",x"6d",x"49",x"6d",x"b2",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"45",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"6e",x"45",x"45",x"49",x"49",x"92",x"49",x"49",x"b6",x"92",x"b6",x"49",x"49",x"b2",x"49",x"92",x"49",x"92",x"69",x"49",x"b6",x"db",x"49",x"49",x"b6",x"8d",x"92",x"49",x"6d",x"49",x"b2",x"b6",x"49",x"69",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"45",x"6d",x"24",x"6d",x"49",x"92",x"6e",x"49",x"6d",x"49",x"92",x"92",x"49",x"49",x"b6",x"b6",x"69",x"92",x"49",x"49",x"db",x"b6",x"69",x"49",x"b2",x"49",x"6d",x"49",x"b6",x"49",x"49",x"b7",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"69",x"49",x"25",x"24",x"24",x"92",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"45",x"25",x"25",x"24",x"25",x"25",x"49",x"6e",x"69",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"45",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"6d",x"49",x"6d",x"24",x"49",x"92",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"b6",x"92",x"92",x"49",x"8d",x"b6",x"b6",x"49",x"69",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"b6",x"b6",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"92",x"45",x"49",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"6d",x"49",x"49",x"45",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"45",x"69",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"92",x"49",x"92",x"b6",x"69",x"49",x"b6",x"b6",x"6d",x"69",x"6d",x"49",x"b6",x"92",x"6d",x"49",x"92",x"92",x"92",x"49",x"49",x"6d",x"49",x"6d",x"69",x"b6",x"49",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"45",x"69",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"45",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"72",x"6d",x"49",x"49",x"69",x"b6",x"49",x"45",x"25",x"49",x"24",x"45",x"24",x"49",x"6d",x"49",x"24",x"24",x"49",x"6e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"24",x"49",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"92",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"6d",x"92",x"b6",x"49",x"49",x"92",x"49",x"92",x"49",x"92",x"6d",x"6d",x"92",x"b6",x"69",x"69",x"b6",x"b6",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"24",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"49",x"69",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"92",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"69",x"6d",x"49",x"49",x"8e",x"92",x"49",x"92",x"49",x"b6",x"92",x"6d",x"49",x"db",x"b6",x"6d",x"6d",x"92",x"49",x"6d",x"69",x"b6",x"49",x"49",x"b6",x"b6",x"49",x"49",x"6d",x"69",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"92",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"25",x"45",x"49",x"b6",x"49",x"45",x"25",x"49",x"24",x"45",x"24",x"49",x"6d",x"49",x"24",x"24",x"25",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"24",x"49",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"69",x"49",x"49",x"25",x"25",x"49",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"92",x"49",x"49",x"92",x"92",x"b6",x"69",x"6d",x"b6",x"db",x"49",x"69",x"b2",x"b6",x"49",x"6d",x"69",x"92",x"69",x"49",x"49",x"92",x"6e",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"24",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"45",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"49",x"49",x"45",x"8e",x"6d",x"6d",x"8e",x"92",x"49",x"8e",x"49",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"45",x"24",x"24",x"49",x"49",x"24",x"49",x"8e",x"49",x"6d",x"49",x"92",x"92",x"49",x"92",x"8e",x"b6",x"49",x"92",x"49",x"b6",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"49",x"92",x"92",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"b2",x"49",x"49",x"b6",x"6d",x"b6",x"49",x"49",x"92",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"49",x"b6",x"49",x"25",x"45",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"24",x"49",x"45",x"49",x"6d",x"24",x"24",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"db",x"92",x"92",x"49",x"49",x"b6",x"b2",x"6d",x"49",x"92",x"6d",x"92",x"49",x"b6",x"6d",x"92",x"69",x"b2",x"6d",x"6d",x"92",x"92",x"49",x"92",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"69",x"24",x"49",x"6d",x"49",x"92",x"49",x"69",x"24",x"6d",x"24",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"25",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"49",x"92",x"69",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"45",x"49",x"49",x"24",x"6d",x"49",x"49",x"69",x"49",x"6d",x"92",x"49",x"92",x"92",x"b6",x"69",x"b2",x"6d",x"b6",x"6d",x"92",x"49",x"6d",x"6d",x"b6",x"49",x"69",x"db",x"db",x"49",x"49",x"b6",x"6d",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"24",x"6d",x"49",x"8e",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"25",x"b2",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"45",x"b6",x"49",x"25",x"49",x"49",x"25",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"25",x"49",x"49",x"24",x"49",x"49",x"49",x"92",x"49",x"25",x"44",x"49",x"b6",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"6e",x"49",x"6d",x"49",x"49",x"6e",x"49",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"69",x"6d",x"92",x"b6",x"49",x"6d",x"b2",x"db",x"49",x"6d",x"92",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"92",x"45",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"45",x"45",x"6d",x"6d",x"49",x"92",x"45",x"92",x"6d",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"24",x"69",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"45",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"25",x"24",x"49",x"69",x"6d",x"49",x"92",x"49",x"92",x"92",x"49",x"6d",x"6d",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"92",x"6d",x"b2",x"92",x"92",x"69",x"b6",x"92",x"b6",x"6d",x"92",x"6d",x"8d",x"6d",x"6d",x"49",x"49",x"92",x"69",x"92",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"92",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"45",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"25",x"49",x"49",x"25",x"25",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"8e"),
     (x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"92",x"fb",x"69",x"45",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"49",x"25",x"45",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"69",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"69",x"24",x"24",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"b6",x"92",x"db",x"69",x"49",x"db",x"b6",x"6d",x"6d",x"b2",x"b2",x"b6",x"49",x"6d",x"92",x"b2",x"69",x"92",x"6d",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"45",x"49",x"6d",x"6d",x"8e",x"49",x"6d",x"92",x"6d",x"24",x"6d",x"49",x"49",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"25",x"49",x"45",x"6d",x"6d",x"6d",x"49",x"8e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"25",x"6d",x"6d",x"49",x"92",x"92",x"49",x"49",x"6e",x"92",x"49",x"92",x"69",x"92",x"6d",x"92",x"49",x"b6",x"92",x"b6",x"6d",x"6d",x"b6",x"db",x"49",x"6d",x"b6",x"6d",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"25",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"25",x"49",x"49",x"45",x"25",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"6d",x"69",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"d7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"6d",x"25",x"49",x"25",x"25",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"49",x"69",x"6d",x"49",x"92",x"6d",x"b2",x"49",x"8d",x"6d",x"92",x"69",x"92",x"49",x"92",x"49",x"69",x"49",x"92",x"49",x"6d",x"49",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"45",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"92",x"b6",x"49",x"6d",x"92",x"92",x"69",x"92",x"6d",x"8d",x"6d",x"92",x"49",x"92",x"6d",x"92",x"49",x"49",x"92",x"92",x"6d",x"49",x"92",x"92",x"b6",x"49",x"49",x"92",x"6e",x"b6",x"49",x"49",x"6d",x"49",x"92",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"29",x"24",x"24",x"92",x"6d",x"45",x"45",x"49",x"45",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"92",x"6d",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"6d",x"49",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"49",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"6d",x"49",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"b6",x"92",x"8e",x"49",x"6d",x"92",x"b7",x"69",x"6d",x"b6",x"92",x"b6",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"49",x"92",x"92",x"92",x"49",x"92",x"b2",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"45",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"92",x"92",x"6d",x"69",x"49",x"49",x"6d",x"69",x"49",x"25",x"24",x"25",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"db",x"b2",x"69",x"92",x"b6",x"b6",x"6d",x"92",x"92",x"b6",x"6d",x"92",x"b6",x"b6",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"92",x"49",x"49",x"44",x"45",x"25",x"49",x"6d",x"24",x"25",x"25",x"24",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"92",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"6d",x"6d",x"6d",x"92",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"49",x"45",x"25",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"92",x"49",x"49",x"b6",x"6d",x"6d",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"49",x"92",x"92",x"b6",x"49",x"92",x"92",x"6d",x"49",x"92",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"25",x"49",x"45",x"49",x"92",x"6d",x"92",x"49",x"92",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"25",x"24",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"45",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"69",x"24",x"6d",x"25",x"25",x"49",x"24",x"6d",x"49",x"49",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"6d",x"49",x"6d",x"6d",x"92",x"6d",x"6e",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"25",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"49",x"49",x"49",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"92",x"69",x"92",x"92",x"b6",x"6d",x"b6",x"92",x"b6",x"6d",x"49",x"b6",x"b6",x"69",x"49",x"b6",x"92",x"b6",x"49",x"49",x"b6",x"92",x"6d",x"49",x"49",x"b6",x"6d",x"6d",x"49",x"49",x"92",x"49",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"b6",x"49",x"49",x"24",x"49",x"25",x"49",x"6d",x"24",x"49",x"49",x"24",x"25",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"6d",x"92",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"45",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"92",x"6d",x"b6",x"49",x"49",x"b2",x"6d",x"92",x"69",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"92",x"49",x"92",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"25",x"6e",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"92",x"92",x"8e",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"8d",x"6d",x"6d",x"69",x"49",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"b6",x"49",x"49",x"45",x"49",x"25",x"6d",x"6d",x"24",x"49",x"49",x"25",x"24",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92"),
     (x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"db",x"6d",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"25",x"25",x"45",x"24",x"49",x"db",x"49",x"25",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"20",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"25",x"49",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"49",x"6d",x"b2",x"b6",x"49",x"49",x"b6",x"b6",x"b6",x"6d",x"6d",x"92",x"b6",x"69",x"6d",x"92",x"92",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"92",x"49",x"69",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"6d",x"49",x"92",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"25",x"25",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"45",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"49",x"49",x"6d",x"92",x"6d",x"49",x"8e",x"49",x"49",x"49",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"b6",x"49",x"6d",x"92",x"b6",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"b6",x"db",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"92",x"6d",x"b6",x"49",x"49",x"6d",x"49",x"92",x"49",x"45",x"25",x"6d",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"db",x"6d",x"49",x"45",x"49",x"45",x"6d",x"49",x"24",x"45",x"49",x"49",x"25",x"45",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"92"),
     (x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b7",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"25",x"49",x"45",x"24",x"49",x"db",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"69",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"25",x"49",x"49",x"92",x"6d",x"6e",x"49",x"49",x"92",x"6d",x"b6",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"92",x"69",x"69",x"b6",x"b6",x"6d",x"6d",x"92",x"b6",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"49",x"49",x"6d",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"20",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"49",x"49",x"6d",x"92",x"92",x"49",x"92",x"49",x"6d",x"49",x"25",x"49",x"49",x"49",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"49",x"24",x"6d",x"92",x"49",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"69",x"92",x"49",x"92",x"b6",x"49",x"69",x"b6",x"b6",x"6d",x"92",x"92",x"92",x"6d",x"92",x"92",x"b6",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"92",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"24",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"25",x"49",x"49",x"25",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"92"),
     (x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"25",x"25",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"45",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"25",x"24",x"25",x"6d",x"45",x"49",x"49",x"49",x"6e",x"49",x"6d",x"49",x"49",x"92",x"92",x"b6",x"49",x"49",x"b6",x"92",x"92",x"6d",x"91",x"92",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"b6",x"49",x"6d",x"92",x"b6",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"6d",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"25",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"92",x"92",x"49",x"b6",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"92",x"b2",x"49",x"49",x"b6",x"92",x"92",x"49",x"49",x"b6",x"92",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"6d",x"49",x"92",x"24",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"25",x"24",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"25",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"db",x"b6",x"6d",x"49",x"69",x"6d",x"b6",x"92"),
     (x"b6",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"92",x"49",x"92",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"49",x"92",x"69",x"49",x"6d",x"49",x"92",x"92",x"b6",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"92",x"92",x"49",x"92",x"49",x"92",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"b6",x"49",x"92",x"49",x"8e",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"6d",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"6d",x"6e",x"69",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"6d",x"49",x"49",x"b6",x"92",x"49",x"92",x"6d",x"8e",x"6d",x"92",x"6d",x"b2",x"92",x"b6",x"6d",x"92",x"b6",x"db",x"6d",x"49",x"b6",x"b6",x"6d",x"49",x"6d",x"49",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"25",x"25",x"49",x"8e",x"24",x"24",x"24",x"49",x"24",x"25",x"25",x"6e",x"b6",x"69",x"49",x"49",x"69",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"d7",x"6d",x"69",x"6d",x"8e",x"b6",x"92"),
     (x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"db",x"92",x"92",x"69",x"8e",x"49",x"b6",x"6d",x"92",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"b6",x"b6",x"49",x"8e",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"49",x"45",x"6d",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"49",x"8e",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"25",x"6d",x"6d",x"49",x"25",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"49",x"24",x"6d",x"6d",x"49",x"6d",x"49",x"69",x"92",x"49",x"6d",x"92",x"b6",x"49",x"b6",x"b6",x"8e",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"49",x"8e",x"6d",x"6d",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"b6",x"6d",x"b6",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"00",x"20",x"20",x"00",x"20",x"00",x"24",x"24",x"00",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"49",x"25",x"49",x"49",x"92",x"24",x"24",x"49",x"49",x"25",x"45",x"25",x"6d",x"b6",x"92",x"6d",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"92",x"db",x"92"),
     (x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"20",x"20",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"49",x"25",x"25",x"92",x"6d",x"92",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"b6",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"8d",x"49",x"b6",x"b6",x"6d",x"49",x"92",x"b6",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"49",x"24",x"6d",x"69",x"49",x"6d",x"6d",x"69",x"6d",x"49",x"6d",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"8e",x"b6",x"49",x"b6",x"92",x"6d",x"49",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"92",x"db",x"49",x"49",x"b6",x"b2",x"8e",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"69",x"92",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"b6",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"b6",x"db",x"92"),
     (x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"49",x"45",x"24",x"25",x"49",x"25",x"45",x"49",x"49",x"44",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"6d",x"49",x"6d",x"25",x"49",x"49",x"25",x"92",x"49",x"49",x"6d",x"49",x"49",x"b6",x"b6",x"49",x"49",x"6d",x"49",x"92",x"6d",x"92",x"49",x"49",x"db",x"b6",x"6d",x"49",x"92",x"49",x"92",x"92",x"49",x"49",x"92",x"92",x"49",x"92",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"24",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"92",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"b6",x"6d",x"6d",x"b6",x"b6",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"25",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"92",x"92",x"6e",x"92",x"92",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"92",x"92",x"b7",x"fb",x"92"),
     (x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"49",x"49",x"24",x"24",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"20",x"00",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"6d",x"24",x"24",x"25",x"24",x"24",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"92",x"49",x"69",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"49",x"b6",x"49",x"92",x"92",x"49",x"49",x"6e",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"25",x"49",x"49",x"24",x"45",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"6d",x"24",x"8e",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"45",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"25",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"6d",x"49",x"24",x"6e",x"49",x"6d",x"8e",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"b6",x"b6",x"49",x"49",x"b6",x"6d",x"92",x"49",x"92",x"6d",x"92",x"92",x"b6",x"49",x"49",x"92",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"29",x"24",x"24",x"25",x"6d",x"b6",x"25",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"6e",x"6d",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"b6",x"b6",x"db",x"ff",x"92"),
     (x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"25",x"49",x"49",x"25",x"24",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"25",x"25",x"24",x"25",x"6d",x"24",x"45",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"92",x"b6",x"49",x"49",x"92",x"49",x"92",x"49",x"92",x"49",x"49",x"b6",x"92",x"92",x"6d",x"92",x"49",x"92",x"92",x"b6",x"49",x"92",x"49",x"6d",x"b6",x"49",x"49",x"92",x"49",x"49",x"6d",x"25",x"49",x"25",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"24",x"49",x"6d",x"49",x"92",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"6d",x"24",x"49",x"24",x"25",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"45",x"24",x"49",x"49",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"b6",x"b6",x"49",x"49",x"6d",x"6d",x"92",x"92",x"49",x"6d",x"db",x"92",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"b6",x"92",x"6d",x"49",x"45",x"49",x"49",x"92",x"24",x"24",x"24",x"25",x"24",x"8e",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"00",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"db",x"db",x"b7",x"db",x"ff",x"92"),
     (x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"44",x"49",x"49",x"49",x"db",x"49",x"45",x"49",x"49",x"25",x"24",x"25",x"92",x"25",x"25",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"25",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"92",x"49",x"49",x"b6",x"92",x"6e",x"49",x"6e",x"49",x"92",x"92",x"92",x"49",x"6d",x"49",x"92",x"92",x"92",x"49",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"6d",x"25",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"49",x"24",x"8e",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"6d",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"b6",x"92",x"49",x"49",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"b6",x"92",x"6d",x"49",x"92",x"49",x"6d",x"92",x"b6",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"25",x"49",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"20",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"25",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"96",x"b6",x"b6",x"b6",x"db",x"ff",x"92"),
     (x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"25",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"45",x"25",x"25",x"92",x"49",x"25",x"25",x"49",x"b2",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"6d",x"45",x"25",x"49",x"25",x"25",x"92",x"49",x"6d",x"49",x"49",x"92",x"6d",x"92",x"49",x"6d",x"49",x"49",x"b6",x"92",x"92",x"69",x"6e",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"49",x"69",x"92",x"92",x"49",x"92",x"49",x"6e",x"92",x"49",x"6d",x"49",x"49",x"6d",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"b6",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"49",x"45",x"6e",x"49",x"49",x"92",x"49",x"92",x"6d",x"49",x"92",x"49",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"49",x"49",x"db",x"92",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"6e",x"49",x"49",x"6d",x"49",x"92",x"25",x"24",x"25",x"45",x"45",x"92",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"45",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"6d",x"db",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"92"),
     (x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"25",x"49",x"49",x"49",x"92",x"db",x"49",x"45",x"49",x"49",x"49",x"25",x"24",x"92",x"49",x"49",x"49",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"6e",x"25",x"49",x"49",x"49",x"69",x"6e",x"92",x"49",x"49",x"6d",x"49",x"49",x"db",x"92",x"6d",x"49",x"92",x"49",x"6d",x"b6",x"b6",x"6d",x"6d",x"49",x"49",x"b6",x"b7",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"6d",x"92",x"25",x"49",x"49",x"24",x"49",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"6d",x"49",x"6d",x"6d",x"b6",x"49",x"92",x"6d",x"92",x"6d",x"92",x"49",x"49",x"b6",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"45",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"92"),
     (x"25",x"24",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"b7",x"45",x"49",x"45",x"49",x"25",x"24",x"24",x"92",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"6d",x"49",x"49",x"db",x"b6",x"6d",x"6d",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"45",x"25",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"49",x"92",x"49",x"49",x"b6",x"92",x"92",x"49",x"49",x"49",x"49",x"92",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"49",x"24",x"24",x"24",x"49",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"ff",x"92"),
     (x"49",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"b6",x"b6",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"92",x"6d",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"20",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"6d",x"24",x"24",x"45",x"24",x"24",x"92",x"6d",x"6d",x"49",x"49",x"69",x"49",x"49",x"b6",x"92",x"6d",x"49",x"6d",x"49",x"49",x"db",x"b6",x"6d",x"49",x"6d",x"49",x"92",x"92",x"92",x"49",x"6d",x"49",x"92",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"92",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"25",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6e",x"49",x"6e",x"92",x"49",x"49",x"92",x"6d",x"92",x"6d",x"92",x"49",x"6d",x"6d",x"8e",x"6d",x"49",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"24",x"25",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"d7",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"92"),
     (x"49",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"92",x"db",x"b2",x"45",x"49",x"49",x"25",x"25",x"25",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"25",x"25",x"49",x"25",x"49",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"92",x"49",x"92",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"45",x"45",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"92",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"69",x"8e",x"49",x"92",x"49",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"6d",x"db",x"92"),
     (x"49",x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"6d",x"6d",x"b6",x"db",x"92",x"25",x"49",x"49",x"25",x"25",x"25",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"6d",x"49",x"25",x"49",x"25",x"49",x"6d",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6e",x"49",x"6d",x"49",x"6d",x"92",x"92",x"6d",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"25",x"6d",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"25",x"45",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"49",x"24",x"44",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"25",x"6d",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"25",x"6d",x"24",x"49",x"49",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"92",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"92",x"92",x"49",x"8e",x"49",x"49",x"92",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"25",x"25",x"24",x"49",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"b6",x"6d",x"49",x"49",x"45",x"49",x"49",x"45",x"6d",x"6d",x"49",x"25",x"45",x"49",x"6d",x"db",x"6d"),
     (x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"92",x"6d",x"6d",x"92",x"92",x"92",x"25",x"25",x"45",x"25",x"24",x"25",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"6d",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"6d",x"45",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"b6",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6e",x"b2",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"45",x"6d",x"69",x"6d",x"24",x"6d",x"24",x"25",x"6d",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"25",x"49",x"24",x"24",x"6d",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6e",x"24",x"49",x"24",x"25",x"25",x"24",x"49",x"6d",x"24",x"24",x"49",x"49",x"49",x"69",x"49",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"69",x"45",x"6d",x"24",x"6d",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"45",x"49",x"45",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6e",x"6d",x"92",x"6d",x"92",x"49",x"49",x"92",x"49",x"92",x"6d",x"b6",x"49",x"49",x"69",x"49",x"6d",x"6d",x"92",x"49",x"45",x"24",x"49",x"49",x"6d",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"b6",x"6d",x"49",x"49",x"45",x"49",x"49",x"25",x"6d",x"49",x"25",x"25",x"25",x"49",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6e",x"b2",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"25",x"25",x"24",x"24",x"25",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"25",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"25",x"49",x"45",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"69",x"45",x"49",x"6d",x"24",x"92",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"6d",x"6d",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"92",x"49",x"24",x"49",x"24",x"24",x"45",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"92",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"49",x"6d",x"6e",x"6d",x"49",x"92",x"24",x"6d",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"25",x"49",x"49",x"25",x"49",x"49",x"92",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"b6",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"20",x"20",x"24",x"8e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"48",x"45",x"49",x"49",x"45",x"45",x"6d",x"49",x"24",x"25",x"25",x"25",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"6d",x"92",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"25",x"24",x"25",x"25",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"69",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"6e",x"49",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"49",x"6d",x"8e",x"92",x"49",x"6d",x"24",x"6d",x"25",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"6d",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"25",x"45",x"49",x"b6",x"49",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"45",x"24",x"69",x"24",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"6e",x"6d",x"b6",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"8d",x"48",x"45",x"49",x"49",x"25",x"49",x"6d",x"25",x"24",x"25",x"25",x"25",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"92",x"92",x"6d",x"69",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"b7",x"49",x"25",x"24",x"25",x"49",x"49",x"25",x"25",x"24",x"25",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"92",x"6e",x"49",x"6d",x"49",x"49",x"6e",x"49",x"92",x"92",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"45",x"49",x"25",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"49",x"92",x"6e",x"6d",x"92",x"49",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"25",x"6d",x"25",x"25",x"25",x"25",x"24",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"25",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"92",x"49",x"44",x"49",x"49",x"25",x"49",x"6d",x"24",x"49",x"25",x"25",x"24",x"49",x"d7",x"6d"),
     (x"49",x"49",x"49",x"92",x"b6",x"8e",x"6d",x"6d",x"d7",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"25",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"45",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"69",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"25",x"25",x"24",x"45",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"92",x"92",x"49",x"6d",x"69",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"25",x"24",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"6d",x"49",x"24",x"24",x"49",x"49",x"45",x"25",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"49",x"25",x"49",x"25",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"6d",x"49",x"45",x"49",x"6d",x"49",x"24",x"24",x"25",x"24",x"45",x"25",x"b2",x"92",x"49",x"45",x"49",x"49",x"25",x"6d",x"49",x"24",x"49",x"25",x"25",x"24",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"8e",x"d7",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"45",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"20",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6e",x"6d",x"6d",x"92",x"6d",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6e",x"6d",x"6d",x"49",x"6d",x"49",x"8e",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"69",x"49",x"92",x"6d",x"92",x"92",x"6d",x"49",x"6d",x"45",x"49",x"49",x"45",x"49",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"25",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6e",x"6d",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"49",x"49",x"6e",x"25",x"24",x"24",x"45",x"25",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"92",x"49",x"92",x"45",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"b6",x"b6",x"6d",x"b6",x"92",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"b6",x"24",x"6d",x"49",x"25",x"24",x"49",x"6d",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"92",x"6d",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"25",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"92",x"25",x"24",x"24",x"49",x"49",x"49",x"25",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"49",x"49",x"25",x"25",x"49",x"d6",x"8d"),
     (x"49",x"69",x"49",x"6d",x"db",x"b6",x"92",x"92",x"b6",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"49",x"49",x"d7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"25",x"24",x"49",x"25",x"49",x"49",x"24",x"49",x"b6",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"8e",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"24",x"69",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"6d",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"49",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"24",x"6d",x"25",x"25",x"24",x"25",x"24",x"49",x"49",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"25",x"24",x"24",x"49",x"49",x"49",x"45",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"45",x"49",x"49",x"49",x"25",x"49",x"db",x"91"),
     (x"49",x"69",x"49",x"6d",x"db",x"db",x"92",x"92",x"b6",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"b7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6e",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"6d",x"25",x"24",x"49",x"25",x"25",x"49",x"49",x"49",x"92",x"49",x"6e",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6e",x"49",x"6e",x"6e",x"49",x"92",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"24",x"6d",x"49",x"49",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"6d",x"24",x"6d",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"6e",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"6d",x"25",x"6d",x"49",x"25",x"25",x"25",x"45",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"6d",x"92",x"25",x"24",x"24",x"49",x"49",x"49",x"45",x"92",x"db",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"91"),
     (x"49",x"49",x"49",x"6d",x"db",x"db",x"96",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"45",x"49",x"24",x"24",x"6d",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6e",x"20",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"92",x"92",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"45",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"92",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"25",x"6d",x"92",x"25",x"24",x"24",x"49",x"49",x"49",x"45",x"6e",x"db",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"92"),
     (x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"25",x"6e",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"6e",x"69",x"49",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"6d",x"b6",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"6d",x"25",x"49",x"49",x"92",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"29",x"24",x"25",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"6d",x"69",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"da",x"92"),
     (x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"25",x"49",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"49",x"92",x"b2",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"20",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"25",x"49",x"24",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"25",x"6d",x"25",x"49",x"6d",x"49",x"6d",x"24",x"49",x"24",x"6d",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"20",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"24",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"45",x"25",x"49",x"49",x"25",x"6d",x"49",x"92",x"49",x"49",x"6e",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"20",x"00",x"24",x"20",x"00",x"00",x"20",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"8e",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6"),
     (x"49",x"49",x"49",x"49",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"25",x"49",x"25",x"24",x"49",x"49",x"92",x"49",x"49",x"6d",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"6d",x"25",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"92",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"69",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"45",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"25",x"45",x"6d",x"6d",x"6d",x"6d",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"45",x"6e",x"49",x"49",x"6e",x"49",x"69",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6e",x"49",x"92",x"49",x"49",x"49",x"25",x"24",x"25",x"25",x"24",x"49",x"24",x"49",x"6d",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6e",x"6e",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"6d",x"6e",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6"),
     (x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"45",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"49",x"49",x"25",x"24",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"25",x"6d",x"49",x"49",x"6d",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"25",x"20",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"24",x"49",x"25",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"69",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"49",x"6e",x"6d",x"25",x"49",x"49",x"49",x"25",x"49",x"45",x"49",x"49",x"49",x"6d",x"49",x"6d",x"69",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"69",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6"),
     (x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"25",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"25",x"25",x"49",x"45",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"25",x"6d",x"92",x"25",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"24",x"45",x"25",x"45",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6d",x"69",x"6d",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"49",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"69",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"49",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"29",x"24",x"49",x"25",x"25",x"6e",x"49",x"92",x"6d",x"49",x"6d",x"6d",x"24",x"6d",x"49",x"25",x"49",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"6d",x"6d",x"92",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"25",x"25",x"49",x"45",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"d7"),
     (x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"92",x"92",x"49",x"25",x"25",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"49",x"45",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"6d",x"49",x"25",x"49",x"25",x"24",x"49",x"49",x"25",x"25",x"49",x"25",x"24",x"45",x"49",x"24",x"25",x"6d",x"24",x"49",x"6e",x"25",x"92",x"69",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"6d",x"6d",x"69",x"49",x"92",x"25",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"25",x"24",x"24",x"49",x"49",x"6d",x"49",x"d7",x"49",x"24",x"24",x"49",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"6d",x"6e",x"6d",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"6e",x"b2",x"6d",x"24",x"49",x"24",x"49",x"49",x"25",x"24",x"45",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"6d",x"49",x"49",x"6d",x"24",x"49",x"25",x"25",x"49",x"25",x"49",x"24",x"24",x"25",x"24",x"49",x"45",x"25",x"49",x"49",x"6d",x"69",x"6e",x"49",x"49",x"92",x"25",x"24",x"24",x"24",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"24",x"24",x"24",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"45",x"45",x"45",x"49",x"25",x"45",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"92",x"b6",x"24",x"24",x"49",x"49",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"92",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"24",x"49",x"25",x"45",x"24",x"25",x"45",x"25",x"24",x"24",x"24",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"6d",x"6d",x"8e",x"49",x"49",x"b6",x"45",x"49",x"b6",x"6d",x"49",x"92",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"6d",x"24",x"49",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"6d",x"45",x"6d",x"6d",x"92",x"49",x"49",x"49",x"69",x"6d",x"45",x"49",x"45",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"6d",x"49",x"49",x"6e",x"49",x"24",x"92",x"24",x"24",x"49",x"49",x"25",x"45",x"49",x"24",x"24",x"49",x"24",x"25",x"49",x"6d",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"25",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"25",x"6d",x"49",x"25",x"24",x"45",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"25",x"49",x"49",x"49",x"25",x"6d",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"25",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"8e",x"6d",x"49",x"92",x"b6",x"25",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"6d",x"49",x"6d",x"24",x"24",x"25",x"24",x"25",x"49",x"92",x"b2",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"6d",x"8e",x"6d",x"69",x"49",x"45",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"45",x"6d",x"b2",x"b6",x"45",x"69",x"49",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"24",x"6e",x"24",x"6d",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"25",x"49",x"49",x"25",x"49",x"24",x"49",x"25",x"49",x"49",x"69",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"00",x"20",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"49",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"25",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"6d",x"24",x"6d",x"24",x"49",x"25",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"24",x"49",x"49",x"6d",x"49",x"49",x"24",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"6e",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"24",x"49",x"45",x"24",x"49",x"24",x"24",x"25",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"24",x"92",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"6d",x"49",x"25",x"8e",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"25",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"25",x"49",x"6d",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"6e",x"49",x"49",x"45",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"d7",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"49",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"6e",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"b6",x"92",x"6d",x"b6",x"24",x"49",x"6d",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"25",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"24",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"45",x"45",x"45",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"fb",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"b6",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"04",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"49",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"49",x"6e",x"24",x"49",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"92",x"6d",x"92",x"92",x"49",x"25",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"8e",x"45",x"49",x"49",x"49",x"49",x"92",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"45",x"45",x"24",x"49",x"6d",x"25",x"25",x"24",x"24",x"24",x"25",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff"),
     (x"49",x"49",x"49",x"49",x"49",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"29",x"92",x"6d",x"6d",x"49",x"6d",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"b7",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"49",x"00",x"20",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"49",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"45",x"69",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"b6",x"24",x"49",x"49",x"8e",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"6d",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"00",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"6e",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"44",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"6d",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"49",x"24",x"6d",x"49",x"24",x"6d",x"24",x"6d",x"6d",x"24",x"6e",x"25",x"49",x"6e",x"49",x"49",x"6d",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b7",x"b7"),
     (x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"92",x"b6",x"92",x"6d",x"29",x"49",x"49",x"49",x"45",x"44",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"6d",x"49",x"24",x"6d",x"6d",x"24",x"49",x"6d",x"24",x"49",x"6d",x"45",x"49",x"49",x"45",x"6d",x"49",x"49",x"49",x"24",x"6d",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"92",x"6d",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"20",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"69",x"49",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"d7",x"49",x"49",x"49",x"49",x"6e",x"49",x"24",x"49",x"25",x"24",x"24",x"25",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"92",x"92",x"92",x"6e",x"6d",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"20",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"49",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"25",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"6d",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"b6",x"49",x"49",x"49",x"49",x"92",x"45",x"24",x"25",x"25",x"25",x"25",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"6d",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"6e",x"49",x"49",x"6e",x"24",x"45",x"6d",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"49",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"49",x"25",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"25",x"25",x"25",x"25",x"49",x"25",x"49",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"b6",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"69",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"49",x"24",x"00",x"25",x"49",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"49",x"49",x"24",x"6d",x"49",x"45",x"6d",x"24",x"45",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"20",x"25",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"25",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"20",x"00",x"00",x"00",x"49",x"25",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6e",x"6d",x"6d",x"92",x"6d",x"45",x"25",x"25",x"24",x"49",x"25",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"4d",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"24",x"49",x"49",x"25",x"25",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"45",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"20",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"25",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"49",x"45",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"25",x"24",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"6d",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"69",x"6d",x"92",x"6e",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"45",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"20",x"00",x"00",x"00",x"25",x"25",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6e",x"6d",x"6e",x"b6",x"49",x"49",x"45",x"25",x"25",x"49",x"25",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"45",x"45",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"25",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"69",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"69",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"69",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"69",x"24",x"49",x"24",x"49",x"24",x"45",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"24",x"6d",x"49",x"24",x"6d",x"49",x"24",x"49",x"6d",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"45",x"25",x"49",x"25",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"44",x"49",x"24",x"25",x"45",x"49",x"b6",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"24",x"24",x"45",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"24",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"45",x"49",x"24",x"6d",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"49",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"69",x"24",x"24",x"49",x"25",x"24",x"49",x"69",x"24",x"49",x"24",x"49",x"49",x"45",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"24",x"29",x"4d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"45",x"49",x"25",x"45",x"49",x"49",x"b6",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"25",x"45",x"00",x"00",x"49",x"24",x"00",x"24",x"49",x"24",x"00",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"45",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"49",x"45",x"24",x"69",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"24",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"49",x"b6",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"69",x"49",x"49",x"49",x"49",x"25",x"49",x"69",x"24",x"49",x"24",x"49",x"24",x"6d",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"20",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"24",x"24",x"24"),
     (x"49",x"49",x"49",x"69",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"24",x"25",x"45",x"24",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"25",x"49",x"24",x"49",x"25",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"00",x"20",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"25",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"69",x"25",x"6d",x"49",x"6d",x"49",x"24",x"6d",x"49",x"6d",x"25",x"24",x"49",x"24",x"49",x"24",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"45",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"6d",x"49",x"24",x"6d",x"49",x"6d",x"24",x"69",x"69",x"49",x"49",x"24",x"69",x"49",x"6d",x"6d",x"24",x"45",x"24",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"00",x"24",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24"),
     (x"6d",x"6d",x"49",x"69",x"8d",x"ff",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"6d",x"45",x"49",x"49",x"6d",x"db",x"6e",x"25",x"25",x"49",x"24",x"49",x"25",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"24",x"20",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"24",x"49",x"24",x"6d",x"6d",x"24",x"6d",x"45",x"6d",x"69",x"24",x"49",x"49",x"6d",x"24",x"49",x"6d",x"25",x"6d",x"49",x"49",x"25",x"49",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"db",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"25",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"45",x"6d",x"24",x"6d",x"6d",x"45",x"45",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"45",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"20",x"49",x"49",x"24",x"24",x"6d",x"20",x"00",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"49",x"24"),
     (x"6d",x"6d",x"69",x"6d",x"91",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"72",x"25",x"25",x"25",x"24",x"25",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"45",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"6d",x"6d",x"25",x"6d",x"45",x"49",x"6d",x"45",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"92",x"49",x"24",x"6d",x"49",x"24",x"45",x"24",x"24",x"25",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"45",x"25",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"6d",x"49",x"49",x"6d",x"45",x"6d",x"49",x"49",x"6d",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"45",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"24",x"24"),
     (x"92",x"6d",x"6d",x"6d",x"8d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"49",x"49",x"49",x"25",x"6d",x"6d",x"49",x"49",x"6e",x"92",x"72",x"49",x"25",x"25",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"00",x"24",x"49",x"24",x"00",x"49",x"49",x"00",x"24",x"49",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"24",x"45",x"24",x"6d",x"49",x"49",x"49",x"24",x"45",x"69",x"6d",x"45",x"6d",x"45",x"6d",x"6e",x"45",x"69",x"49",x"6d",x"45",x"92",x"6d",x"49",x"49",x"69",x"45",x"49",x"25",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"45",x"25",x"49",x"6d",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"6d",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"69",x"92",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"69",x"6d",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"45",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"24",x"24"),
     (x"b6",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"69",x"49",x"6e",x"6d",x"6d",x"49",x"24",x"24",x"49",x"25",x"24",x"49",x"b6",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"45",x"00",x"00",x"25",x"45",x"00",x"00",x"49",x"24",x"00",x"24",x"49",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"24",x"69",x"24",x"69",x"49",x"24",x"49",x"45",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"25",x"49",x"49",x"25",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"6d",x"92",x"49",x"49",x"92",x"92",x"6d",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"45",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"69",x"6d",x"45",x"8e",x"6d",x"49",x"69",x"24",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"00",x"20",x"24",x"45",x"00",x"24",x"49",x"24",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"92",x"49",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"24",x"24"),
     (x"db",x"92",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"24",x"49",x"45",x"24",x"49",x"b6",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"24",x"49",x"24",x"6d",x"6d",x"25",x"49",x"49",x"6d",x"69",x"69",x"49",x"92",x"92",x"49",x"92",x"69",x"49",x"6d",x"6d",x"49",x"49",x"8e",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"24",x"25",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"b6",x"6d",x"6d",x"69",x"92",x"49",x"6d",x"49",x"45",x"25",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"25",x"6d",x"6d",x"6d",x"8e",x"6d",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"8e",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"45",x"6d",x"49",x"49",x"6d",x"24",x"45",x"24",x"49",x"45",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"45",x"00",x"00",x"49",x"24",x"00",x"24",x"49",x"00",x"00",x"45",x"49",x"00",x"24",x"49",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"6e",x"6e",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"69",x"49",x"69",x"92",x"6d",x"49",x"49",x"49",x"24",x"24"),
     (x"db",x"b6",x"92",x"92",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"49",x"49",x"45",x"49",x"25",x"b6",x"6e",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"25",x"44",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"00",x"20",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"6d",x"6d",x"45",x"49",x"49",x"92",x"92",x"49",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"45",x"49",x"49",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"b6",x"49",x"49",x"24",x"24",x"45",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"92",x"6d",x"49",x"6d",x"49",x"8e",x"6d",x"45",x"49",x"45",x"49",x"49",x"69",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"20",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"24"),
     (x"b6",x"db",x"b2",x"b6",x"db",x"ff",x"db",x"b6",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"25",x"49",x"49",x"b6",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"49",x"00",x"20",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"25",x"45",x"24",x"6d",x"6d",x"24",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"b2",x"8e",x"49",x"8e",x"6d",x"49",x"6d",x"49",x"49",x"6e",x"6d",x"69",x"92",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"49",x"45",x"49",x"49",x"92",x"49",x"92",x"92",x"6d",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"8e",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6e",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"8d",x"92",x"49",x"6d",x"8e",x"6d",x"6d",x"45",x"6d",x"6e",x"25",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"20",x"49",x"25",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"24",x"24",x"00",x"20",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"04",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"45",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"6d",x"6e",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"24"),
     (x"92",x"fb",x"d7",x"db",x"db",x"db",x"b6",x"b6",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"49",x"b6",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"20",x"45",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"6d",x"69",x"24",x"25",x"49",x"49",x"6d",x"69",x"49",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"92",x"6d",x"6d",x"69",x"92",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"92",x"b6",x"b6",x"6d",x"49",x"45",x"49",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"b6",x"49",x"69",x"92",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"69",x"49",x"92",x"92",x"49",x"b6",x"92",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"45",x"6d",x"6d",x"25",x"6d",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"25",x"20",x"20",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"25",x"24",x"00",x"49",x"25",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"20",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"49",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"b6",x"92",x"92",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"25",x"24"),
     (x"6d",x"ff",x"db",x"db",x"db",x"b6",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"25",x"49",x"45",x"49",x"49",x"db",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"49",x"b6",x"92",x"24",x"25",x"45",x"24",x"24",x"24",x"25",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"24",x"20",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"6d",x"69",x"45",x"25",x"6d",x"45",x"6d",x"8e",x"49",x"69",x"8e",x"92",x"49",x"92",x"92",x"49",x"49",x"6d",x"69",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"6d",x"49",x"69",x"d7",x"b6",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"92",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"49",x"25",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"24",x"49",x"69",x"49",x"25",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"49",x"92",x"8e",x"49",x"8e",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"69",x"49",x"b2",x"6d",x"49",x"49",x"45",x"49",x"49",x"6d",x"24",x"25",x"24",x"25",x"25",x"45",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"49",x"24",x"00",x"24",x"49",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"6d",x"24",x"20",x"00",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"b6",x"92",x"92",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"25",x"24"),
     (x"6d",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"45",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"20",x"24",x"24",x"24",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"49",x"20",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"6d",x"25",x"69",x"6d",x"45",x"49",x"92",x"92",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"92",x"8e",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"25",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"6d",x"49",x"45",x"92",x"49",x"49",x"49",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6e",x"6d",x"49",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"45",x"49",x"25",x"25",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"92",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"25",x"6d",x"24",x"49",x"24",x"6d",x"45",x"49",x"6d",x"24",x"49",x"6d",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"69",x"49",x"49",x"6d",x"6d",x"6e",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"92",x"b6",x"49",x"6d",x"b6",x"49",x"6d",x"49",x"8e",x"69",x"49",x"45",x"6d",x"6d",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"20",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"92",x"92",x"92",x"d7",x"db",x"6d",x"49",x"49",x"49",x"49",x"25",x"24"),
     (x"6d",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"92",x"6e",x"49",x"24",x"49",x"24",x"49",x"49",x"25",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"25",x"49",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"49",x"69",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"45",x"92",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"6d",x"25",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"25",x"24",x"49",x"49",x"45",x"49",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"45",x"45",x"49",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"25",x"49",x"49",x"6d",x"49",x"49",x"6d",x"69",x"6d",x"49",x"92",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"b6",x"49",x"92",x"6e",x"49",x"b6",x"92",x"49",x"6d",x"92",x"92",x"49",x"6d",x"49",x"49",x"6d",x"45",x"49",x"49",x"6d",x"24",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"20",x"24",x"49",x"20",x"24",x"25",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"45",x"24",x"25",x"25",x"25",x"b6",x"6d",x"48",x"49",x"49",x"49",x"49",x"49",x"6e",x"6d",x"69",x"6d",x"92",x"b6",x"d7",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"24"),
     (x"6d",x"92",x"ff",x"db",x"6e",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"25",x"24",x"24",x"25",x"6e",x"49",x"49",x"6d",x"92",x"49",x"49",x"24",x"49",x"25",x"25",x"49",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"45",x"8e",x"6d",x"49",x"49",x"92",x"6d",x"49",x"92",x"49",x"92",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"92",x"49",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"25",x"49",x"49",x"49",x"49",x"45",x"6d",x"49",x"69",x"49",x"92",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"45",x"24",x"6d",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"92",x"49",x"69",x"92",x"92",x"69",x"92",x"92",x"49",x"92",x"92",x"6d",x"49",x"92",x"b6",x"49",x"b2",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"24",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"00",x"20",x"24",x"20",x"20",x"49",x"25",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"49",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"00",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"25",x"24",x"45",x"25",x"25",x"24",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6e",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"44",x"49",x"24"),
     (x"6d",x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"25",x"24",x"24",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"24",x"25",x"24",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"25",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"25",x"20",x"20",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"6d",x"69",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"49",x"6d",x"b6",x"49",x"92",x"92",x"49",x"92",x"6e",x"6d",x"6d",x"6d",x"92",x"8e",x"6e",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"25",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"8e",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"24",x"92",x"25",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"45",x"25",x"49",x"49",x"6d",x"45",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"49",x"49",x"92",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"49",x"92",x"92",x"69",x"92",x"6d",x"92",x"92",x"69",x"92",x"92",x"49",x"b6",x"92",x"49",x"b6",x"92",x"69",x"49",x"8e",x"92",x"49",x"49",x"45",x"49",x"24",x"69",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"24",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"49",x"24",x"00",x"24",x"25",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"25",x"25",x"25",x"45",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"25",x"49",x"24"),
     (x"6d",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"49",x"49",x"45",x"24",x"49",x"b2",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"92",x"6e",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"6d",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"20",x"00",x"24",x"20",x"20",x"45",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"6d",x"49",x"69",x"24",x"49",x"45",x"6d",x"49",x"8e",x"49",x"8e",x"8e",x"49",x"6d",x"92",x"6d",x"49",x"92",x"8d",x"6d",x"b6",x"49",x"b6",x"92",x"49",x"92",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"92",x"49",x"6d",x"8e",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"24",x"49",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"45",x"45",x"49",x"6d",x"24",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"25",x"45",x"24",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"69",x"6d",x"6d",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"49",x"92",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"6d",x"92",x"6d",x"92",x"6d",x"92",x"92",x"49",x"92",x"b6",x"49",x"b6",x"92",x"49",x"92",x"92",x"8e",x"49",x"b6",x"8e",x"49",x"49",x"6d",x"8e",x"45",x"49",x"25",x"45",x"24",x"69",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"45",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b7",x"49",x"49",x"25",x"25",x"25",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"25",x"45",x"24"),
     (x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"25",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"92",x"b6",x"49",x"6d",x"92",x"8e",x"49",x"6d",x"92",x"92",x"92",x"69",x"92",x"92",x"69",x"6d",x"92",x"92",x"49",x"92",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"69",x"49",x"6d",x"6d",x"6d",x"69",x"6d",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"6e",x"6d",x"49",x"6d",x"92",x"49",x"db",x"6d",x"92",x"6d",x"b2",x"49",x"49",x"6d",x"6d",x"25",x"49",x"6d",x"49",x"49",x"25",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"92",x"6d",x"b6",x"92",x"92",x"6d",x"92",x"b6",x"6d",x"b6",x"92",x"6d",x"6d",x"92",x"8d",x"49",x"b6",x"92",x"49",x"49",x"8e",x"92",x"49",x"8e",x"69",x"6d",x"45",x"69",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"49",x"49",x"45",x"24",x"49",x"49",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"45",x"49",x"6e",x"49",x"25",x"49",x"45",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"24"),
     (x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"45",x"49",x"49",x"49",x"25",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"49",x"6d",x"45",x"49",x"6d",x"8e",x"49",x"92",x"92",x"92",x"49",x"92",x"db",x"49",x"92",x"6d",x"92",x"6d",x"69",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"6d",x"b6",x"6d",x"6d",x"6d",x"92",x"49",x"8e",x"69",x"6d",x"49",x"49",x"6d",x"6d",x"24",x"49",x"25",x"49",x"24",x"24",x"25",x"24",x"25",x"25",x"24",x"49",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"6d",x"69",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"69",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"92",x"49",x"92",x"49",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"92",x"6d",x"92",x"49",x"92",x"8e",x"49",x"69",x"92",x"92",x"6d",x"69",x"92",x"92",x"49",x"92",x"b2",x"49",x"6d",x"6d",x"8d",x"49",x"6d",x"6d",x"69",x"45",x"6d",x"69",x"49",x"24",x"49",x"45",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"20",x"24",x"25",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"25",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"49",x"25",x"24",x"49",x"49",x"25",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"44",x"49",x"45",x"24"),
     (x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"8e",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"25",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"25",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"49",x"6d",x"24",x"45",x"6d",x"6d",x"45",x"49",x"92",x"92",x"49",x"92",x"92",x"92",x"49",x"92",x"d7",x"49",x"92",x"69",x"92",x"b6",x"49",x"b6",x"92",x"92",x"b6",x"49",x"92",x"8d",x"92",x"49",x"92",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"b2",x"92",x"b2",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"b2",x"6d",x"49",x"25",x"45",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"b6",x"92",x"69",x"92",x"8e",x"92",x"69",x"8e",x"6d",x"69",x"69",x"6d",x"49",x"49",x"49",x"24",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"49",x"92",x"8e",x"6d",x"6d",x"6e",x"6d",x"92",x"b6",x"6d",x"92",x"92",x"6d",x"92",x"69",x"92",x"b6",x"49",x"92",x"92",x"69",x"6e",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"8e",x"49",x"49",x"24",x"6d",x"6d",x"49",x"24",x"49",x"45",x"24",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"44",x"49",x"45",x"49"),
     (x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"25",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"69",x"49",x"25",x"49",x"6d",x"6d",x"49",x"49",x"8e",x"92",x"49",x"92",x"92",x"92",x"49",x"b2",x"b2",x"69",x"b6",x"49",x"b6",x"b6",x"6d",x"b6",x"69",x"b2",x"8e",x"6d",x"49",x"92",x"6d",x"92",x"6d",x"6e",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"6d",x"49",x"69",x"6d",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"24",x"25",x"24",x"45",x"24",x"49",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"45",x"24",x"49",x"69",x"49",x"6d",x"49",x"6d",x"6d",x"b6",x"49",x"6d",x"49",x"24",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"20",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"92",x"49",x"49",x"6d",x"24",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"92",x"92",x"6d",x"92",x"6d",x"49",x"92",x"92",x"6d",x"6d",x"49",x"b2",x"b6",x"69",x"b6",x"92",x"6d",x"8e",x"49",x"6d",x"49",x"92",x"49",x"6d",x"69",x"49",x"49",x"6d",x"49",x"25",x"25",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"25",x"49",x"49",x"25",x"49",x"92",x"b7",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"d7",x"92",x"49",x"49",x"49",x"45",x"45",x"49",x"45",x"49"),
     (x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"92",x"db",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"45",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"8e",x"92",x"49",x"92",x"92",x"b6",x"6d",x"92",x"6d",x"92",x"92",x"6d",x"b6",x"92",x"92",x"b2",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"6d",x"49",x"49",x"6d",x"6d",x"69",x"6d",x"92",x"6d",x"49",x"92",x"6d",x"92",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"45",x"24",x"49",x"49",x"24",x"6d",x"25",x"6d",x"92",x"6d",x"92",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"8e",x"49",x"92",x"49",x"6d",x"6d",x"49",x"49",x"8e",x"69",x"6d",x"49",x"24",x"49",x"45",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"b6",x"6d",x"92",x"49",x"92",x"92",x"92",x"92",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"92",x"49",x"49",x"92",x"92",x"49",x"45",x"6d",x"6d",x"24",x"24",x"49",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"69",x"24",x"45",x"49",x"45",x"49",x"25",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"44",x"49",x"49",x"45",x"49"),
     (x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"69",x"6d",x"92",x"db",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"92",x"92",x"49",x"6d",x"92",x"92",x"49",x"6d",x"69",x"92",x"8e",x"6d",x"6d",x"6d",x"92",x"6d",x"92",x"49",x"92",x"49",x"92",x"6d",x"6e",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"25",x"24",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"92",x"6d",x"92",x"6d",x"b6",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"6d",x"49",x"49",x"45",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"b6",x"6d",x"92",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"92",x"49",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"92",x"6d",x"49",x"92",x"6d",x"49",x"92",x"49",x"92",x"b6",x"49",x"49",x"92",x"92",x"49",x"49",x"6d",x"8e",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"6d",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"25",x"6d"),
     (x"49",x"49",x"49",x"92",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"92",x"b2",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"6e",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"45",x"24",x"6d",x"49",x"6d",x"25",x"6d",x"6d",x"6d",x"49",x"8e",x"8e",x"6d",x"49",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"6d",x"8d",x"6d",x"6d",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6e",x"49",x"6d",x"49",x"49",x"49",x"49",x"25",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"49",x"49",x"92",x"8e",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"45",x"49",x"24",x"25",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"25",x"49",x"45",x"49",x"24",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"92",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"69",x"24",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"49",x"92",x"92",x"92",x"b6",x"49",x"b2",x"6d",x"b6",x"6d",x"69",x"6d",x"6d",x"b6",x"92",x"49",x"92",x"49",x"92",x"b6",x"49",x"69",x"92",x"92",x"49",x"6d",x"49",x"6d",x"45",x"49",x"49",x"49",x"24",x"45",x"49",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"24",x"24",x"24",x"00",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"44",x"49",x"45",x"49",x"49",x"49",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"49",x"49",x"49",x"6d",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b2",x"b2",x"b2",x"92",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"24",x"00",x"20",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"24",x"6d",x"49",x"6d",x"45",x"49",x"92",x"92",x"49",x"49",x"92",x"6d",x"49",x"92",x"49",x"8e",x"92",x"49",x"6d",x"49",x"92",x"6d",x"92",x"92",x"49",x"92",x"49",x"92",x"b6",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"6d",x"49",x"69",x"49",x"49",x"69",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"8e",x"6d",x"49",x"49",x"49",x"24",x"45",x"49",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"45",x"24",x"25",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"69",x"8e",x"6d",x"6d",x"49",x"92",x"6d",x"69",x"49",x"49",x"6d",x"45",x"6d",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"49",x"6d",x"49",x"92",x"92",x"6d",x"92",x"49",x"b2",x"92",x"92",x"92",x"49",x"92",x"6d",x"92",x"92",x"49",x"6e",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"45",x"69",x"25",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"24",x"24",x"24",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"49",x"45",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"92",x"6e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"49",x"49",x"45",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"24",x"25",x"24",x"24",x"24",x"45",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"20",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"b2",x"92",x"6d",x"92",x"49",x"92",x"92",x"92",x"b6",x"49",x"6d",x"49",x"92",x"92",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"69",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"69",x"49",x"92",x"49",x"49",x"45",x"49",x"69",x"25",x"24",x"49",x"45",x"49",x"24",x"25",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"25",x"6d",x"49",x"49",x"92",x"49",x"6d",x"49",x"92",x"6d",x"92",x"49",x"92",x"49",x"92",x"92",x"49",x"92",x"49",x"92",x"92",x"49",x"6d",x"49",x"92",x"92",x"6d",x"49",x"92",x"49",x"6d",x"49",x"49",x"45",x"6d",x"6d",x"45",x"24",x"49",x"49",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"45",x"45",x"24",x"24",x"24",x"24",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"6d",x"b6",x"49",x"24",x"24",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db"),
     (x"49",x"49",x"45",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"45",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"00",x"24",x"24",x"6d",x"00",x"00",x"00",x"24",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"69",x"49",x"45",x"6d",x"49",x"6d",x"49",x"69",x"49",x"6d",x"6d",x"6d",x"49",x"92",x"49",x"b6",x"b6",x"49",x"6d",x"49",x"92",x"b2",x"6d",x"b6",x"49",x"92",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"49",x"45",x"49",x"6d",x"45",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"45",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"45",x"25",x"49",x"24",x"24",x"24",x"45",x"25",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"92",x"6d",x"24",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"49",x"92",x"49",x"92",x"6d",x"92",x"b6",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"92",x"45",x"24",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"00",x"69",x"24",x"24",x"24",x"20",x"20",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"b6",x"49",x"24",x"24",x"25",x"29",x"49",x"49",x"49",x"25",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db"),
     (x"49",x"49",x"44",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b7",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6e",x"92",x"6d",x"b6",x"49",x"6e",x"49",x"6d",x"6d",x"92",x"92",x"49",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"25",x"69",x"49",x"24",x"49",x"49",x"24",x"49",x"25",x"25",x"24",x"49",x"49",x"49",x"69",x"49",x"25",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"69",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"45",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"45",x"6d",x"25",x"92",x"24",x"49",x"92",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"b6",x"6d",x"92",x"6e",x"49",x"6d",x"49",x"b6",x"92",x"92",x"92",x"49",x"49",x"8d",x"6d",x"49",x"49",x"49",x"6d",x"6e",x"8e",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"6d",x"24",x"24",x"24",x"20",x"20",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"49",x"24",x"25",x"25",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff"),
     (x"48",x"49",x"44",x"49",x"92",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"25",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"24",x"24",x"49",x"25",x"69",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"20",x"00",x"00",x"49",x"00",x"00",x"00",x"24",x"20",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"6d",x"6d",x"45",x"49",x"92",x"69",x"6d",x"92",x"49",x"49",x"92",x"6d",x"6d",x"92",x"49",x"92",x"49",x"6d",x"92",x"6d",x"92",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"24",x"69",x"49",x"69",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"49",x"24",x"24",x"25",x"45",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"6d",x"24",x"6d",x"49",x"92",x"24",x"49",x"49",x"45",x"49",x"69",x"24",x"49",x"6d",x"49",x"49",x"24",x"49",x"45",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"6d",x"25",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"92",x"49",x"92",x"49",x"b6",x"6d",x"92",x"92",x"49",x"92",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"25",x"69",x"49",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"20",x"00",x"24",x"20",x"6d",x"20",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"92",x"b6",x"49",x"49",x"45",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff"),
     (x"24",x"48",x"49",x"49",x"6d",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"6e",x"49",x"25",x"49",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"b6",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"69",x"00",x"00",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"92",x"92",x"6d",x"b6",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"92",x"6d",x"92",x"49",x"6d",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"49",x"49",x"6d",x"49",x"45",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"25",x"49",x"25",x"49",x"49",x"49",x"6d",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"92",x"49",x"92",x"92",x"49",x"45",x"6d",x"6d",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff"),
     (x"24",x"44",x"49",x"49",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"25",x"49",x"45",x"25",x"49",x"6d",x"49",x"49",x"49",x"92",x"db",x"b6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"24",x"49",x"24",x"49",x"45",x"49",x"45",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"69",x"49",x"49",x"24",x"49",x"24",x"49",x"92",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6e",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"45",x"24",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"25",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"6d",x"69",x"49",x"45",x"49",x"25",x"49",x"6d",x"6d",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"20",x"00",x"24",x"25",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"d7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff"),
     (x"48",x"24",x"49",x"49",x"49",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"24",x"49",x"45",x"49",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"6d",x"25",x"45",x"25",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"b6",x"92",x"69",x"92",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"45",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"24",x"25",x"49",x"49",x"24",x"45",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"92",x"49",x"6d",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6e",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"92",x"92",x"69",x"25",x"49",x"49",x"6d",x"6d",x"69",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"db"),
     (x"49",x"24",x"48",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"24",x"24",x"49",x"44",x"49",x"6d",x"6d",x"24",x"25",x"25",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"20",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"6d",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"6e",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"25",x"6d",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"25",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"25",x"49",x"45",x"6d",x"49",x"49",x"25",x"49",x"49",x"49",x"6d",x"49",x"92",x"49",x"6e",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6d",x"69",x"25",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db"),
     (x"49",x"44",x"48",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"72",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"25",x"49",x"45",x"24",x"45",x"6d",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"45",x"24",x"49",x"49",x"49",x"24",x"24",x"6d",x"49",x"6d",x"6d",x"24",x"49",x"49",x"49",x"6d",x"49",x"92",x"92",x"49",x"92",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"45",x"24",x"49",x"24",x"49",x"24",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"45",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"45",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"92",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"24",x"49",x"24",x"49",x"49",x"6d",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"6d",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"b7"),
     (x"49",x"49",x"48",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"92",x"25",x"49",x"49",x"45",x"24",x"45",x"49",x"db",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"49",x"24",x"49",x"6d",x"49",x"25",x"49",x"24",x"69",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"25",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"6d",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"92",x"49",x"6e",x"6d",x"69",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"6d",x"45",x"6d",x"49",x"24",x"6d",x"45",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"b6",x"b7",x"96",x"b6"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"8e",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"25",x"49",x"49",x"24",x"49",x"69",x"b7",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"49",x"24",x"25",x"49",x"45",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"24",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"49",x"69",x"49",x"69",x"49",x"6e",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"45",x"69",x"6d",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"24",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"6d",x"b2",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"69",x"49",x"69",x"49",x"49",x"49",x"6d",x"db",x"92",x"92",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"b6",x"6d",x"49",x"24",x"24",x"25",x"49",x"49",x"49",x"45",x"49",x"6d",x"b6",x"6e",x"49",x"24",x"45",x"45",x"24",x"49",x"49",x"b7",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"6d",x"49",x"49",x"6d",x"25",x"49",x"24",x"49",x"24",x"25",x"49",x"25",x"49",x"25",x"6d",x"24",x"6d",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"6d",x"49",x"6e",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"b7",x"49",x"24",x"25",x"24",x"25",x"49",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6e",x"6e",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"25",x"24",x"25",x"25",x"24",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"44",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"25",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"45",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"49",x"25",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"6d",x"25",x"49",x"25",x"6d",x"6d",x"49",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"b6",x"49",x"24",x"25",x"24",x"49",x"49",x"24",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"25",x"24",x"25",x"45",x"24",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"44",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"b6",x"24",x"24",x"25",x"24",x"49",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"24",x"20",x"45",x"25",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"20",x"20",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"45",x"49",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"6d",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"25",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"49",x"25",x"49",x"49",x"24",x"6d",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6e",x"45",x"24",x"24",x"25",x"49",x"49",x"25",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"92",x"69",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"4d",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"25",x"24",x"24",x"49",x"49",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"d7",x"49",x"24",x"25",x"24",x"49",x"25",x"45",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"00",x"24",x"24",x"24",x"6d",x"00",x"24",x"20",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"49",x"24",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"49",x"45",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"20",x"20",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"25",x"24",x"25",x"25",x"25",x"24",x"25",x"24",x"49",x"24",x"92",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"25",x"24",x"25",x"24",x"24",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"20",x"20",x"20",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b7",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"24",x"24",x"49",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"92",x"6e",x"49",x"24",x"24",x"24",x"49",x"24",x"45",x"b2",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"69",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"6d",x"92",x"92",x"6d",x"92",x"6d",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"25",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"69",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"20",x"00",x"00",x"49",x"24",x"24",x"20",x"20",x"20",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"4d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"45",x"45",x"49",x"24",x"24",x"92",x"92",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"20",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"92",x"6d",x"6d",x"92",x"92",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"24",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"24",x"24",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"29",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"6d",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d"),
     (x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"45",x"25",x"44",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"25",x"24",x"49",x"49",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"04",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"8e",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"49",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d"),
     (x"92",x"49",x"49",x"49",x"69",x"6d",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"49",x"45",x"24",x"24",x"44",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"20",x"20",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"6e",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"25",x"24",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"24",x"24",x"00",x"00",x"24",x"49",x"00",x"24",x"24",x"20",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"d7",x"8d",x"6d",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"25",x"6d"),
     (x"92",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"45",x"49",x"49",x"44",x"24",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"92",x"49",x"6d",x"6d",x"92",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"db",x"b6",x"8d",x"6d",x"69",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"29",x"6d"),
     (x"92",x"92",x"49",x"6d",x"69",x"6d",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"49",x"45",x"24",x"24",x"49",x"49",x"db",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"69",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"92",x"49",x"6d",x"92",x"6d",x"8d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"6d",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"20",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"db",x"b6",x"92",x"8e",x"6d",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"29",x"92"),
     (x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"8d",x"d6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"49",x"49",x"24",x"24",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"45",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"8d",x"69",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"b7",x"b6",x"92",x"92",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"49",x"92",x"92",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"92",x"49",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"25",x"25",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"6d",x"6d",x"49",x"6d",x"8e",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"20",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6e",x"b6",x"b7",x"b2",x"b6",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db"),
     (x"49",x"6d",x"b2",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"45",x"00",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"92",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"49",x"b6",x"92",x"92",x"92",x"49",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"69",x"49",x"6d",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"b7",x"b6",x"b7",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db"),
     (x"49",x"6d",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"20",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"20",x"49",x"00",x"24",x"00",x"00",x"24",x"24",x"49",x"00",x"20",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"45",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"45",x"45",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6e",x"49",x"92",x"6d",x"6d",x"92",x"b2",x"6d",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"25",x"24",x"49",x"24",x"49",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"20",x"25",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"49",x"49",x"24",x"24",x"45",x"25",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"4d",x"49",x"92",x"b7",x"db",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db"),
     (x"49",x"49",x"6e",x"b6",x"92",x"6d",x"92",x"92",x"db",x"db",x"db",x"92",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"45",x"49",x"44",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"00",x"24",x"20",x"6d",x"00",x"20",x"00",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"25",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"49",x"6d",x"92",x"6d",x"92",x"49",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"92",x"49",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"45",x"20",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"48",x"24",x"24",x"24",x"45",x"24",x"24",x"92",x"6d",x"49",x"45",x"24",x"25",x"49",x"25",x"49",x"db",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"4d",x"49",x"49",x"6e",x"b6",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6"),
     (x"49",x"49",x"6d",x"b6",x"b2",x"6d",x"92",x"92",x"b7",x"db",x"b6",x"b6",x"6d",x"49",x"6d",x"6d",x"69",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"45",x"49",x"45",x"49",x"49",x"24",x"92",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"00",x"00",x"24",x"24",x"45",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"49",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"b2",x"49",x"b2",x"6d",x"92",x"6d",x"92",x"92",x"49",x"69",x"92",x"69",x"49",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"49",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"b6",x"49",x"49",x"25",x"25",x"25",x"49",x"25",x"49",x"db",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92"),
     (x"49",x"49",x"49",x"92",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"92",x"b6",x"92",x"49",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"45",x"49",x"45",x"6d",x"92",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"45",x"6d",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"8e",x"6d",x"49",x"b6",x"92",x"49",x"6d",x"6d",x"92",x"6d",x"69",x"92",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"00",x"45",x"00",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"20",x"20",x"24",x"20",x"24",x"24",x"6d",x"24",x"24",x"24",x"00",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"24",x"49",x"49",x"45",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d"),
     (x"49",x"49",x"49",x"6d",x"b6",x"b6",x"b6",x"b6",x"b6",x"b6",x"72",x"92",x"92",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"20",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"92",x"6d",x"6d",x"49",x"b6",x"92",x"49",x"8e",x"92",x"6d",x"49",x"92",x"6d",x"49",x"92",x"45",x"6d",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"45",x"45",x"20",x"24",x"24",x"20",x"20",x"49",x"45",x"24",x"24",x"24",x"24",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8e",x"92",x"db",x"92",x"49",x"69",x"6d",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"49"),
     (x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"b7",x"b6",x"96",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"24",x"24",x"24",x"49",x"48",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"6d",x"69",x"25",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"8e",x"69",x"6d",x"92",x"49",x"8d",x"6d",x"49",x"6d",x"92",x"69",x"6d",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"20",x"00",x"00",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"48",x"24",x"25",x"45",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6e",x"b6",x"92",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"db",x"b6",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"92",x"49",x"8e",x"49",x"49",x"6d",x"92",x"49",x"92",x"92",x"49",x"6d",x"92",x"49",x"92",x"49",x"92",x"49",x"6d",x"6d",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"25",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"44",x"25",x"45",x"45",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"92",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"b6",x"92",x"4d",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"db",x"db",x"8e",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"6d",x"49",x"49",x"6e",x"49",x"6d",x"6d",x"49",x"49",x"92",x"6d",x"49",x"92",x"6d",x"69",x"92",x"49",x"92",x"8e",x"49",x"49",x"6d",x"49",x"49",x"49",x"24",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"49",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"db",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"b7",x"49",x"45",x"24",x"45",x"45",x"49",x"49",x"92",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"8e",x"6d",x"49",x"6d",x"92",x"db",x"db",x"92",x"6d",x"49",x"6d",x"69",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"24",x"49",x"24",x"45",x"6d",x"b6",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"24",x"49",x"45",x"6d",x"6d",x"49",x"8e",x"6d",x"49",x"69",x"92",x"49",x"6d",x"6d",x"49",x"92",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"45",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"49",x"49",x"24",x"45",x"49",x"49",x"4d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6e",x"b7",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"6d",x"8d",x"b7",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"24",x"49",x"25",x"49",x"44",x"45",x"49",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"04",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"25",x"00",x"24",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"25",x"69",x"69",x"49",x"6d",x"49",x"6d",x"92",x"49",x"8e",x"92",x"49",x"6d",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"45",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"8e",x"48",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"6d",x"6e",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"45",x"49",x"49",x"6e",x"b7",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"8d",x"92",x"b6",x"b2",x"6d",x"6e",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"45",x"49",x"24",x"24",x"24",x"49",x"b6",x"6d",x"25",x"24",x"24",x"24",x"24",x"45",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"49",x"24",x"00",x"24",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"6d",x"49",x"6d",x"8e",x"45",x"6d",x"6d",x"49",x"6d",x"6d",x"69",x"69",x"69",x"49",x"6d",x"45",x"69",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"24",x"24",x"24",x"45",x"24",x"25",x"49",x"b6",x"92",x"49",x"24",x"45",x"24",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"25",x"25",x"25",x"49",x"6e",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"69",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"fb",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"25",x"49",x"24",x"24",x"24",x"48",x"8d",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"24",x"24",x"24",x"6d",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"20",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"45",x"69",x"45",x"69",x"69",x"45",x"6d",x"69",x"69",x"49",x"49",x"6d",x"49",x"49",x"6d",x"45",x"49",x"8e",x"45",x"6d",x"24",x"49",x"45",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"20",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"6d",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"25",x"49",x"24",x"25",x"49",x"92",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"d6",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"b6",x"b6",x"b6",x"92",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"69",x"92",x"db",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"d7",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"d7",x"92",x"25",x"25",x"25",x"24",x"25",x"24",x"6d",x"b7",x"49",x"24",x"24",x"24",x"25",x"25",x"49",x"b7",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"20",x"49",x"24",x"00",x"00",x"04",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"25",x"6d",x"49",x"49",x"45",x"49",x"6d",x"45",x"6d",x"6d",x"45",x"6d",x"49",x"69",x"24",x"49",x"45",x"45",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"92",x"6d",x"49",x"25",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"6e",x"6d",x"92",x"6d",x"45",x"45",x"45",x"49",x"25",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"49",x"49"),
     (x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"db",x"b7",x"b6",x"6e",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"69",x"92",x"db",x"92",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"49",x"24",x"24",x"45",x"24",x"44",x"49",x"b7",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"24",x"6d",x"49",x"24",x"6d",x"49",x"69",x"45",x"49",x"92",x"25",x"6d",x"25",x"6d",x"49",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"25",x"24",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"25",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"92",x"49",x"45",x"49",x"45",x"49",x"25",x"49",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49"),
     (x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"b7",x"6d",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"6e",x"49",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"45",x"24",x"25",x"45",x"45",x"25",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"45",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"24",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"24",x"00",x"20",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"25",x"49",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"6d",x"45",x"49",x"49",x"49",x"25",x"25",x"6d",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49"),
     (x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"6e",x"92",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b7",x"6d",x"49",x"49",x"45",x"45",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"24",x"25",x"25",x"24",x"45",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"69",x"6d",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"b6",x"49",x"49",x"49",x"45",x"49",x"25",x"25",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49"),
     (x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"25",x"45",x"49",x"6d",x"b6",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"6e",x"6d",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"45",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"45",x"24",x"49",x"6d",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"20",x"24",x"20",x"00",x"20",x"24",x"49",x"24",x"24",x"20",x"24",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"b2",x"6d",x"49",x"45",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49"),
     (x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6e",x"92",x"49",x"45",x"49",x"49",x"49",x"25",x"49",x"6d",x"92",x"49",x"25",x"49",x"49",x"25",x"25",x"25",x"6d",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"24",x"20",x"25",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"49",x"25",x"49",x"25",x"49",x"45",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"25",x"25",x"24",x"24",x"25",x"6d",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49"),
     (x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"b6",x"92",x"49",x"49",x"49",x"45",x"49",x"6d",x"6d",x"6d",x"92",x"6d",x"45",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"6e",x"24",x"24",x"24",x"49",x"49",x"29",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"49",x"25",x"25",x"25",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"da",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"b7",x"92",x"49",x"25",x"49",x"49",x"45",x"49",x"92",x"92",x"92",x"6d",x"25",x"24",x"24",x"24",x"49",x"6d",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"20",x"20",x"45",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"45",x"24",x"24",x"49",x"25",x"24",x"24",x"45",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"20",x"25",x"20",x"24",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"49",x"25",x"25",x"24",x"24",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"45",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49"),
     (x"b6",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"25",x"49",x"49",x"45",x"45",x"6d",x"b6",x"b2",x"6d",x"25",x"25",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"4d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"20",x"00",x"20",x"20",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"20",x"24",x"69",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"25",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"45",x"49",x"24",x"45",x"49",x"49",x"24",x"45",x"24",x"45",x"24",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"24",x"25",x"25",x"25",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"45",x"49",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"b7",x"6d",x"24",x"25",x"49",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"29",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"25",x"24",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"24",x"49",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"25",x"25",x"49",x"25",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"db",x"6e",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"6d",x"db",x"6e",x"25",x"24",x"25",x"25",x"45",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"45",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"45",x"49",x"25",x"45",x"49",x"45",x"24",x"6d",x"b6",x"49",x"49",x"49",x"45",x"49",x"25",x"45",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"92",x"6e",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"24",x"49",x"49",x"49",x"25",x"25",x"92",x"6e",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"25",x"20",x"24",x"24",x"24",x"49",x"24",x"69",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"20",x"25",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"24",x"00",x"25",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"6d",x"b6",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"44",x"6d",x"db",x"49",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"25",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"20",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"45",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"25",x"00",x"00",x"49",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"45",x"24",x"24",x"25",x"24",x"49",x"b2",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"b6",x"45",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"b6",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"45",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"44",x"49",x"b6",x"6d",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"20",x"49",x"24",x"24",x"24",x"00",x"49",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"44",x"24",x"24",x"24",x"49",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"45",x"49",x"25",x"49",x"49",x"49",x"25",x"92",x"92",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"da",x"6d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"24",x"49",x"49",x"49",x"45",x"49",x"44",x"6d",x"b6",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"25",x"24",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"00",x"24",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"b6",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"45",x"b6",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"45",x"b6",x"49",x"24",x"49",x"25",x"24",x"24",x"45",x"49",x"b6",x"49",x"24",x"45",x"24",x"24",x"24",x"25",x"49",x"92",x"24",x"24",x"25",x"49",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"45",x"20",x"00",x"24",x"00",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"20",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"20",x"25",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"24",x"00",x"20",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"8e",x"49",x"25",x"25",x"45",x"24",x"24",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"ff",x"ff",x"8d",x"69",x"49",x"69",x"49",x"49",x"49",x"b6"),
     (x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"49",x"24",x"49",x"44",x"49",x"b6",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"25",x"49",x"24",x"25",x"24",x"45",x"b6",x"25",x"24",x"25",x"25",x"24",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"00",x"25",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"20",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"20",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"6d",x"24",x"49",x"24",x"24",x"25",x"25",x"25",x"b6",x"49",x"49",x"45",x"49",x"45",x"24",x"24",x"49",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"b6",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db"),
     (x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"24",x"45",x"49",x"45",x"45",x"49",x"49",x"49",x"b6",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"44",x"92",x"49",x"24",x"49",x"49",x"24",x"25",x"25",x"49",x"b6",x"49",x"25",x"25",x"24",x"25",x"49",x"48",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"48",x"24",x"24",x"24",x"25",x"25",x"69",x"b6",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"6d",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"db"),
     (x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"45",x"25",x"49",x"49",x"49",x"6d",x"92",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"6d",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"24",x"24",x"24",x"25",x"49",x"24",x"49",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"49",x"24",x"20",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"b6",x"6d",x"49",x"49",x"45",x"45",x"45",x"25",x"45",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"69",x"49",x"6d",x"49",x"6d",x"b6",x"ff",x"ff",x"b2",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"b6"),
     (x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"45",x"45",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"24",x"45",x"49",x"25",x"49",x"49",x"92",x"6d",x"24",x"25",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"20",x"24",x"49",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"db",x"49",x"44",x"45",x"44",x"45",x"45",x"25",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"92",x"ff",x"8e",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"8e",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"b7",x"92"),
     (x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8e",x"24",x"49",x"49",x"25",x"24",x"49",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"00",x"20",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"8e",x"92",x"49",x"49",x"45",x"45",x"45",x"45",x"25",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"db",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d"),
     (x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"49",x"49",x"24",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"20",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"25",x"49",x"49",x"24",x"49",x"45",x"24",x"49",x"49",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"69",x"49",x"49",x"24",x"49",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"25",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"00",x"24",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"45",x"45",x"25",x"49",x"45",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"69",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"25",x"25",x"49",x"24",x"24",x"49",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"25",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"49",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"25",x"24",x"49",x"6d",x"6d",x"25",x"24",x"24",x"49",x"49",x"49",x"25",x"45",x"25",x"49",x"25",x"24",x"24",x"6d",x"69",x"49",x"25",x"24",x"49",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"49",x"24",x"49",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"04",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"b7",x"49",x"45",x"45",x"49",x"45",x"45",x"45",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"69",x"69",x"49",x"6d",x"db",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d"),
     (x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"44",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"49",x"24",x"24",x"49",x"6d",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"04",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"24",x"20",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6e",x"49",x"49",x"24",x"25",x"49",x"49",x"49",x"25",x"45",x"49",x"24",x"49",x"25",x"25",x"25",x"25",x"49",x"24",x"25",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"49",x"20",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"25",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"b6",x"6d",x"6d",x"49",x"49",x"69",x"49",x"69",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"db",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"49",x"6d"),
     (x"49",x"49",x"49",x"49",x"69",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6e",x"25",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"6d",x"25",x"24",x"25",x"24",x"25",x"49",x"6d",x"29",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"25",x"24",x"24",x"6d",x"6d",x"49",x"49",x"45",x"45",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"6d",x"6d",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"6e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"92",x"db",x"ff",x"d6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"b7",x"db",x"bb",x"db",x"db",x"b6",x"6d",x"8d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"d7",x"92",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"29",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"25",x"6d",x"24",x"25",x"6d",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"25",x"6d",x"6d",x"49",x"49",x"25",x"49",x"24",x"24",x"49",x"6d",x"6d",x"25",x"25",x"49",x"6d",x"6d",x"49",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"20",x"20",x"00",x"6d",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"db",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"b7",x"db",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"b6",x"db",x"db",x"b2",x"92",x"92",x"92",x"b6",x"92",x"6d",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"92",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"b6",x"92",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"00",x"49",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"49",x"24",x"49",x"24",x"25",x"25",x"25",x"24",x"49",x"49",x"49",x"24",x"49",x"6d",x"6d",x"49",x"25",x"49",x"49",x"25",x"49",x"92",x"6d",x"49",x"49",x"25",x"92",x"6d",x"6d",x"45",x"29",x"49",x"6d",x"6e",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"25",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"45",x"6d",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"6d",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"25",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"25",x"25",x"25",x"49",x"92",x"49",x"24",x"24",x"25",x"45",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"6d",x"b6",x"db",x"db",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"92",x"db",x"db",x"db",x"92",x"6d",x"6d",x"6e",x"6d",x"92",x"b7",x"b6",x"92",x"b6",x"db",x"db",x"b2",x"92",x"92",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"fb",x"db",x"49",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"29",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"45",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"8e",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"6d",x"24",x"24",x"24",x"00",x"24",x"00",x"45",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"24",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"45",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"45",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"92",x"b6",x"db",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"b7",x"b6",x"db",x"db",x"6d",x"6d",x"6d",x"8e",x"6e",x"b6",x"b6",x"92",x"92",x"b6",x"b6",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"b6",x"ff",x"92",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6e",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"20",x"00",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"49",x"25",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"6d",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"96",x"db",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"b6",x"b6",x"92",x"db",x"b6",x"6d",x"6d",x"6e",x"6d",x"92",x"b6",x"92",x"6e",x"92",x"b6",x"b7",x"db",x"b6",x"b6",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"6e"),
     (x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"92",x"ff",x"db",x"69",x"6d",x"49",x"49",x"69",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6e",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"45",x"49",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"25",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"49",x"24",x"45",x"92",x"6d",x"49",x"49",x"6e",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"24",x"45",x"49",x"49",x"49",x"25",x"25",x"49",x"45",x"24",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"45",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"6e",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"72",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"92",x"db",x"b6",x"92",x"6d",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"ff",x"ff",x"92",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"8d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"6d",x"49",x"24",x"6d",x"6d",x"49",x"45",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"8e",x"49",x"49",x"49",x"92",x"6d",x"6e",x"49",x"49",x"49",x"69",x"49",x"6d",x"69",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"45",x"69",x"6d",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"6d",x"69",x"49",x"49",x"6d",x"8e",x"6d",x"6d",x"96",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"6d",x"92",x"db",x"b6",x"92",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"fb",x"db",x"92",x"6d",x"49",x"6d",x"49",x"49",x"6d",x"b7"),
     (x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"69",x"8d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"db",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"6d",x"24",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"24",x"49",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"24",x"00",x"00",x"00",x"20",x"00",x"49",x"25",x"24",x"00",x"24",x"24",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"45",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"92",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"92",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"24",x"49",x"6d",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"20",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"69",x"6d",x"72",x"6d",x"49",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"92",x"8e",x"6d",x"6d",x"92",x"db",x"b6",x"b6",x"92",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"db"),
     (x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"92",x"ff",x"d7",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"25",x"25",x"49",x"6d",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"29",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"6d",x"6d",x"49",x"24",x"6d",x"6d",x"24",x"24",x"8e",x"49",x"25",x"6d",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"92",x"6d",x"92",x"49",x"49",x"49",x"b6",x"6d",x"92",x"49",x"6d",x"49",x"92",x"8e",x"6e",x"49",x"49",x"49",x"92",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"6e",x"6d",x"49",x"6d",x"49",x"49",x"25",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b2",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"25",x"25",x"45",x"6d",x"b6",x"92",x"6d",x"6e",x"6e",x"6d",x"49",x"49",x"6d",x"92",x"b6",x"92",x"6d",x"8e",x"b6",x"92",x"6d",x"49",x"6d",x"92",x"db",x"b6",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"92",x"ff"),
     (x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"6d",x"6d",x"69",x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"25",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"25",x"25",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6e",x"49",x"49",x"69",x"6d",x"49",x"6d",x"49",x"49",x"49",x"92",x"6e",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"8e",x"24",x"49",x"6d",x"49",x"24",x"49",x"6d",x"49",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"24",x"25",x"25",x"6d",x"b6",x"92",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"92",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"92",x"db",x"db",x"db",x"db",x"92",x"6d",x"6d",x"4d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff"),
     (x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"b6",x"69",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"25",x"25",x"24",x"00",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"69",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"49",x"24",x"25",x"25",x"49",x"49",x"25",x"92",x"6d",x"49",x"6e",x"92",x"6d",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"92",x"6e",x"6e",x"49",x"49",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"92",x"49",x"49",x"49",x"92",x"49",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6d",x"92",x"49",x"6d",x"6e",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"25",x"25",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"20",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"92",x"49",x"25",x"25",x"25",x"25",x"25",x"6e",x"b6",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"b2",x"b6",x"b6",x"6d",x"49",x"49",x"6d",x"6d",x"b6",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"4d",x"4d",x"49",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"ff",x"ff"),
     (x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"6e",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"25",x"24",x"24",x"24",x"24",x"25",x"25",x"49",x"b6",x"25",x"24",x"24",x"24",x"45",x"45",x"24",x"69",x"b2",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"25",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"24",x"45",x"25",x"6d",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6d",x"92",x"92",x"b6",x"49",x"6d",x"49",x"b6",x"92",x"b6",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"92",x"45",x"49",x"92",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6e",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"6d",x"92",x"6d",x"25",x"25",x"25",x"25",x"24",x"25",x"92",x"b6",x"96",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"b7",x"ff",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"6e",x"b7",x"ff",x"ff",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"4d",x"b6",x"ff",x"db"),
     (x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6e",x"49",x"49",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6e",x"6d",x"49",x"49",x"49",x"49",x"6e",x"92",x"6d",x"49",x"25",x"45",x"49",x"6d",x"6e",x"6e",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6e",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"00",x"00",x"24",x"20",x"00",x"49",x"25",x"24",x"00",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"45",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"92",x"92",x"92",x"92",x"49",x"49",x"69",x"49",x"49",x"49",x"b6",x"92",x"92",x"92",x"49",x"49",x"6d",x"92",x"6e",x"92",x"49",x"49",x"49",x"92",x"92",x"92",x"69",x"49",x"49",x"6d",x"8e",x"49",x"8e",x"6d",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"49",x"92",x"92",x"49",x"25",x"24",x"25",x"25",x"24",x"49",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"b7",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"49",x"6d",x"db",x"ff",x"92"),
     (x"ff",x"db",x"ff",x"b6",x"92",x"6d",x"6e",x"6d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"db",x"92",x"6d",x"4d",x"6d",x"6d",x"49",x"49",x"6e",x"92",x"6d",x"45",x"25",x"25",x"49",x"4d",x"92",x"92",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"b6",x"49",x"24",x"45",x"24",x"24",x"49",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"92",x"69",x"24",x"25",x"92",x"6d",x"24",x"24",x"6d",x"6d",x"49",x"45",x"92",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"b6",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"6e",x"6d",x"92",x"92",x"49",x"49",x"49",x"6e",x"49",x"49",x"92",x"92",x"6d",x"92",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"24",x"49",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"b6",x"49",x"25",x"24",x"25",x"25",x"25",x"24",x"49",x"b6",x"b6",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"6e",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"6d",x"49",x"6d",x"49",x"49",x"92",x"ff",x"db",x"6d"),
     (x"ff",x"db",x"ff",x"db",x"b6",x"6d",x"92",x"6d",x"6d",x"91",x"b6",x"ff",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"db",x"b6",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"92",x"6d",x"49",x"25",x"25",x"24",x"49",x"6d",x"92",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"25",x"24",x"24",x"45",x"49",x"6d",x"b6",x"24",x"25",x"24",x"24",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"45",x"25",x"45",x"6d",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"92",x"92",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"92",x"49",x"49",x"49",x"b6",x"92",x"92",x"92",x"49",x"49",x"8e",x"49",x"6d",x"6d",x"92",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"92",x"92",x"49",x"92",x"92",x"49",x"49",x"92",x"6d",x"24",x"49",x"6e",x"6d",x"24",x"49",x"6d",x"6d",x"25",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"00",x"24",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"25",x"24",x"24",x"49",x"25",x"25",x"25",x"6d",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"b7",x"ff",x"92",x"6d"),
     (x"ff",x"db",x"db",x"ff",x"db",x"92",x"92",x"92",x"8d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b7",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"6e",x"92",x"6d",x"49",x"45",x"49",x"25",x"25",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"b6",x"6d",x"24",x"24",x"24",x"25",x"49",x"25",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"b6",x"6d",x"6d",x"8e",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"b6",x"8e",x"db",x"6d",x"49",x"49",x"6d",x"b6",x"92",x"b6",x"49",x"49",x"49",x"b6",x"92",x"b6",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"92",x"b7",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"49",x"25",x"45",x"24",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"6d"),
     (x"db",x"ff",x"bb",x"db",x"db",x"b6",x"92",x"92",x"92",x"8e",x"92",x"b6",x"ff",x"db",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"db",x"b7",x"b6",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"db",x"92",x"6d",x"72",x"92",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"92",x"6e",x"49",x"29",x"49",x"49",x"49",x"25",x"49",x"b7",x"49",x"24",x"25",x"24",x"24",x"25",x"24",x"25",x"6d",x"92",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"69",x"b6",x"45",x"24",x"24",x"24",x"49",x"44",x"49",x"92",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"49",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"6d",x"92",x"49",x"6d",x"6e",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",x"92",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"92",x"69",x"6d",x"6d",x"b6",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"69",x"49",x"49",x"92",x"6d",x"92",x"b6",x"6d",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b2",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"45",x"24",x"49",x"24",x"24",x"24",x"25",x"b6",x"6d",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"92",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"24",x"6d",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"96",x"ff",x"92",x"6d",x"49"),
     (x"db",x"ff",x"bb",x"b6",x"db",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"db",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"6d",x"6d",x"6e",x"92",x"6d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"b6",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"25",x"24",x"25",x"24",x"24",x"25",x"49",x"25",x"92",x"6d",x"24",x"24",x"25",x"24",x"49",x"49",x"45",x"b6",x"92",x"24",x"25",x"25",x"49",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"45",x"49",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"45",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"92",x"92",x"6d",x"db",x"49",x"49",x"49",x"92",x"69",x"49",x"6d",x"92",x"6d",x"6d",x"92",x"49",x"49",x"49",x"b6",x"6d",x"92",x"92",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"b6",x"92",x"db",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6e",x"92",x"49",x"6d",x"92",x"92",x"49",x"49",x"6d",x"6e",x"49",x"49",x"25",x"6d",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"45",x"49",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"45",x"45",x"49",x"25",x"24",x"24",x"49",x"b6",x"49",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"b6",x"92",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"6d",x"49"),
     (x"b6",x"ff",x"db",x"b6",x"b6",x"db",x"d6",x"92",x"92",x"92",x"92",x"92",x"db",x"ff",x"b6",x"b6",x"db",x"b6",x"8d",x"6d",x"6d",x"6d",x"92",x"ff",x"b6",x"92",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"6d",x"49",x"69",x"6d",x"92",x"92",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"6d",x"24",x"45",x"24",x"24",x"24",x"25",x"49",x"49",x"b6",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"b7",x"49",x"25",x"24",x"49",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"92",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"25",x"24",x"49",x"92",x"49",x"24",x"24",x"6d",x"49",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"92",x"b6",x"6d",x"92",x"92",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"92",x"92",x"92",x"b6",x"49",x"49",x"49",x"92",x"b6",x"92",x"db",x"49",x"49",x"6d",x"92",x"b6",x"92",x"db",x"49",x"49",x"49",x"6e",x"6d",x"49",x"49",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"49",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"20",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"25",x"49",x"25",x"24",x"24",x"25",x"b6",x"6d",x"48",x"45",x"25",x"25",x"24",x"25",x"24",x"49",x"b6",x"49",x"24",x"24",x"25",x"45",x"45",x"25",x"24",x"69",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"6d",x"49",x"49"),
     (x"b6",x"db",x"db",x"b6",x"b6",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"d6",x"ff",x"b6",x"b6",x"b6",x"b6",x"92",x"8d",x"6d",x"91",x"92",x"db",x"b6",x"92",x"6e",x"92",x"b6",x"92",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"49",x"49",x"49",x"92",x"b6",x"b6",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6e",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"49",x"24",x"49",x"25",x"49",x"49",x"92",x"92",x"24",x"49",x"24",x"25",x"49",x"49",x"49",x"92",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"25",x"6d",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"20",x"00",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"92",x"6d",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"b2",x"8d",x"db",x"6d",x"6d",x"49",x"49",x"b6",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"92",x"49",x"6d",x"b6",x"6d",x"69",x"6d",x"b6",x"b6",x"92",x"b7",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"92",x"6d",x"92",x"92",x"6d",x"92",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"24",x"6d",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"24",x"25",x"6d",x"b2",x"49",x"49",x"25",x"25",x"25",x"25",x"24",x"6e",x"b6",x"49",x"48",x"24",x"45",x"49",x"45",x"24",x"24",x"b6",x"6d",x"45",x"24",x"25",x"45",x"45",x"45",x"25",x"24",x"b6",x"6d",x"25",x"25",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"6d",x"49",x"49"),
     (x"b6",x"db",x"ff",x"b6",x"92",x"b6",x"db",x"db",x"92",x"92",x"92",x"92",x"b6",x"ff",x"b7",x"92",x"92",x"b6",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"92",x"6d",x"6d",x"92",x"b6",x"92",x"92",x"92",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"92",x"24",x"49",x"25",x"25",x"49",x"24",x"49",x"49",x"d7",x"49",x"25",x"25",x"25",x"49",x"24",x"49",x"6d",x"b7",x"69",x"49",x"24",x"49",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"20",x"20",x"25",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"25",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"92",x"92",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"92",x"92",x"6d",x"8d",x"92",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"92",x"6d",x"49",x"6d",x"db",x"92",x"b6",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"49",x"49",x"49",x"6e",x"49",x"24",x"25",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"25",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"6d",x"49",x"25",x"24",x"25",x"49",x"25",x"49",x"db",x"6d",x"44",x"24",x"45",x"49",x"49",x"25",x"25",x"6d",x"b6",x"49",x"49",x"45",x"45",x"45",x"49",x"49",x"24",x"6d",x"b6",x"49",x"25",x"49",x"49",x"25",x"49",x"49",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49"),
     (x"b6",x"da",x"ff",x"db",x"92",x"92",x"b6",x"db",x"b6",x"92",x"92",x"92",x"b6",x"fb",x"db",x"92",x"92",x"92",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"49",x"25",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"25",x"25",x"49",x"24",x"24",x"49",x"92",x"6e",x"49",x"49",x"45",x"45",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"49",x"6d",x"6e",x"49",x"24",x"49",x"92",x"92",x"25",x"24",x"49",x"b6",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"92",x"92",x"6d",x"b6",x"92",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"b6",x"92",x"92",x"b6",x"49",x"69",x"69",x"b6",x"b6",x"92",x"db",x"69",x"6d",x"6d",x"6d",x"db",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"49",x"6d",x"6d",x"db",x"92",x"b6",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"24",x"25",x"25",x"25",x"25",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"b6",x"49",x"44",x"24",x"24",x"25",x"45",x"25",x"92",x"b6",x"49",x"49",x"45",x"49",x"49",x"25",x"49",x"49",x"b6",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"45",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"45",x"25",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6e",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"6d",x"49",x"49",x"49"),
     (x"b6",x"d6",x"db",x"db",x"92",x"92",x"92",x"b6",x"db",x"b6",x"92",x"92",x"b6",x"db",x"fb",x"92",x"92",x"6e",x"92",x"b6",x"b6",x"92",x"b6",x"b6",x"db",x"92",x"6d",x"6d",x"69",x"6d",x"b6",x"b6",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"b7",x"6d",x"25",x"49",x"49",x"49",x"24",x"24",x"69",x"92",x"49",x"45",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"20",x"24",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"25",x"25",x"49",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"6d",x"b6",x"92",x"b6",x"db",x"49",x"49",x"6d",x"92",x"92",x"6d",x"92",x"92",x"49",x"6d",x"6d",x"92",x"6d",x"6d",x"b6",x"6d",x"6d",x"69",x"92",x"db",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b7",x"92",x"6d",x"92",x"b6",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"92",x"6d",x"45",x"25",x"49",x"92",x"49",x"24",x"25",x"6d",x"8e",x"49",x"25",x"25",x"6d",x"6d",x"6e",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"25",x"24",x"25",x"25",x"6d",x"92",x"49",x"24",x"24",x"25",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"25",x"49",x"49",x"45",x"25",x"6d",x"b6",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"44",x"45",x"49",x"24",x"69",x"db",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"45",x"49",x"d7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49"),
     (x"b6",x"db",x"db",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"b6",x"92",x"b6",x"d6",x"ff",x"b6",x"92",x"6d",x"92",x"92",x"b7",x"b6",x"b6",x"b6",x"fb",x"b6",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"db",x"db",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"24",x"49",x"49",x"45",x"49",x"49",x"24",x"49",x"92",x"6d",x"24",x"25",x"49",x"49",x"49",x"45",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"49",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"25",x"25",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"b7",x"6d",x"49",x"92",x"92",x"6d",x"92",x"b6",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"b6",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"92",x"b6",x"49",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"45",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"24",x"25",x"25",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"44",x"25",x"45",x"b6",x"92",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"db",x"db",x"ff",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"b6",x"b6",x"b6",x"ff",x"b7",x"8e",x"6d",x"6d",x"92",x"b6",x"db",x"b6",x"db",x"db",x"db",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"96",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"b6",x"49",x"45",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"45",x"49",x"49",x"45",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"6d",x"8e",x"92",x"49",x"25",x"49",x"92",x"6d",x"49",x"49",x"92",x"db",x"6d",x"49",x"8e",x"92",x"92",x"92",x"b6",x"92",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"49",x"69",x"49",x"b6",x"b6",x"92",x"db",x"6d",x"49",x"49",x"6d",x"db",x"b6",x"92",x"db",x"6d",x"6d",x"6d",x"69",x"db",x"92",x"b6",x"db",x"6d",x"69",x"6d",x"92",x"6d",x"6d",x"69",x"92",x"db",x"92",x"b6",x"b6",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"45",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"25",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"48",x"45",x"24",x"6d",x"d7",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"db",x"db",x"db",x"db",x"92",x"92",x"6e",x"92",x"b6",x"db",x"db",x"b6",x"db",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"8e",x"6d",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"96",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"24",x"45",x"49",x"25",x"49",x"49",x"49",x"49",x"92",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"24",x"49",x"49",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6e",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"b6",x"92",x"db",x"6d",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"92",x"6d",x"6d",x"6d",x"6d",x"db",x"92",x"92",x"ff",x"49",x"69",x"49",x"6d",x"6d",x"49",x"49",x"49",x"db",x"92",x"6d",x"8e",x"b2",x"6d",x"92",x"b6",x"b2",x"49",x"49",x"92",x"b6",x"6d",x"25",x"25",x"6d",x"92",x"49",x"24",x"49",x"6d",x"92",x"6d",x"49",x"49",x"25",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"4d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"25",x"b7",x"6d",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"db",x"db",x"db",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"db",x"db",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"49",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b6",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"25",x"25",x"24",x"00",x"00",x"00",x"45",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"20",x"20",x"20",x"00",x"00",x"24",x"24",x"00",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"45",x"25",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"92",x"b6",x"92",x"92",x"db",x"49",x"6d",x"49",x"6d",x"92",x"49",x"49",x"6d",x"b6",x"92",x"92",x"db",x"49",x"49",x"6d",x"49",x"db",x"b6",x"92",x"db",x"6d",x"6d",x"69",x"69",x"92",x"6d",x"6d",x"6d",x"b6",x"92",x"92",x"db",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6d",x"92",x"24",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"20",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"4d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"d6",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"b2",x"49",x"49",x"44",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"48"),
     (x"db",x"ff",x"db",x"db",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"44",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"25",x"49",x"49",x"92",x"92",x"92",x"49",x"24",x"49",x"92",x"92",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"92",x"b6",x"92",x"92",x"b6",x"92",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"6d",x"db",x"b6",x"b6",x"ff",x"49",x"49",x"6d",x"6d",x"b6",x"92",x"6d",x"b6",x"6d",x"6d",x"6d",x"69",x"b7",x"b6",x"92",x"fb",x"6d",x"6d",x"6d",x"69",x"b6",x"6d",x"6d",x"69",x"b6",x"b6",x"92",x"b6",x"b6",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"25",x"49",x"25",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"20",x"24",x"45",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"69",x"45",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"b6",x"69",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"28",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48"),
     (x"b6",x"ff",x"fb",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"ff",x"ff",x"db",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"45",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"49",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"45",x"6d",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"92",x"db",x"92",x"b6",x"db",x"6d",x"49",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"b6",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"69",x"92",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"b6",x"b6",x"49",x"49",x"69",x"6d",x"92",x"49",x"49",x"49",x"db",x"b6",x"92",x"92",x"b6",x"6d",x"6d",x"92",x"db",x"6d",x"49",x"49",x"92",x"92",x"49",x"45",x"49",x"6d",x"92",x"6d",x"25",x"49",x"69",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"25",x"49",x"6e",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"92",x"92",x"49",x"49",x"44",x"48",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24"),
     (x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6e",x"b6",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"ff",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"25",x"45",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"20",x"45",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"49",x"24",x"24",x"24",x"45",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"6d",x"db",x"92",x"b2",x"db",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"6d",x"6d",x"db",x"b6",x"b6",x"fb",x"6d",x"69",x"6d",x"6d",x"db",x"b6",x"b2",x"ff",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"6d",x"6d",x"b6",x"8e",x"69",x"6d",x"db",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"92",x"25",x"25",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"45",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"25",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"49",x"49",x"49",x"44",x"49",x"49",x"49",x"49",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"24"),
     (x"6e",x"b6",x"ff",x"ff",x"ff",x"ff",x"b6",x"6e",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"bb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"25",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"8e",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"20",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"25",x"00",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"6d",x"92",x"6e",x"6d",x"49",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"b2",x"b6",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"92",x"69",x"49",x"49",x"69",x"b2",x"db",x"92",x"b2",x"b6",x"69",x"6d",x"6d",x"6d",x"92",x"49",x"49",x"92",x"92",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"69",x"db",x"92",x"6d",x"8d",x"b6",x"6d",x"6d",x"b6",x"db",x"49",x"49",x"49",x"69",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"24",x"49",x"49",x"25",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"24",x"24",x"24",x"25",x"92",x"49",x"49",x"45",x"25",x"49",x"49",x"6d",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"48",x"48",x"49",x"49",x"49",x"44",x"49",x"db",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"24"),
     (x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"6d",x"25",x"25",x"49",x"45",x"6d",x"92",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"b6",x"b6",x"6d",x"6d",x"6d",x"b2",x"49",x"69",x"6d",x"6d",x"db",x"b6",x"b2",x"db",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"92",x"b6",x"6d",x"69",x"49",x"92",x"6d",x"69",x"69",x"49",x"6d",x"b6",x"49",x"49",x"6d",x"b6",x"92",x"6d",x"b6",x"b6",x"6d",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"92",x"92",x"49",x"45",x"49",x"6d",x"b2",x"6d",x"25",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"45",x"25",x"49",x"49",x"6d",x"8e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"48",x"25",x"49"),
     (x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"92",x"6d",x"49",x"6d",x"49",x"49",x"49",x"69",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"25",x"25",x"24",x"49",x"92",x"49",x"24",x"25",x"24",x"49",x"25",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"24",x"20",x"49",x"25",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"49",x"24",x"45",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"db",x"92",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"b6",x"49",x"49",x"49",x"49",x"b2",x"b6",x"92",x"92",x"db",x"6d",x"6d",x"6d",x"6d",x"b6",x"92",x"6d",x"b6",x"b6",x"6d",x"69",x"6d",x"6d",x"ff",x"b6",x"b2",x"d6",x"92",x"49",x"49",x"49",x"b6",x"49",x"69",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"b2",x"25",x"24",x"25",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"69",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"6d",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"d7",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"69",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"49",x"24",x"8e"),
     (x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"b7",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"25",x"49",x"49",x"24",x"6d",x"92",x"25",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"6e",x"25",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"00",x"24",x"24",x"49",x"69",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"6d",x"49",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"6d",x"b7",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"92",x"b6",x"b6",x"92",x"b6",x"b6",x"49",x"49",x"49",x"b6",x"6d",x"49",x"69",x"49",x"6d",x"b6",x"6d",x"49",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"49",x"6d",x"6d",x"49",x"b6",x"92",x"6d",x"92",x"b6",x"49",x"69",x"49",x"92",x"6d",x"69",x"69",x"49",x"92",x"ff",x"92",x"92",x"db",x"92",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"25",x"45",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"00",x"20",x"24",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"44",x"24",x"45",x"24",x"24",x"24",x"24",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"6e",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b7",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6e",x"25",x"24",x"45",x"25",x"49",x"49",x"49",x"92",x"6e",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"db",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"00",x"24",x"49",x"00",x"00",x"24",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"49",x"25",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"ff",x"6d",x"6d",x"6d",x"69",x"6d",x"db",x"92",x"92",x"db",x"6d",x"69",x"6d",x"6d",x"6d",x"ff",x"b6",x"b6",x"ff",x"6d",x"69",x"6d",x"49",x"92",x"6d",x"69",x"49",x"69",x"92",x"db",x"92",x"92",x"92",x"b6",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"45",x"6d",x"6d",x"45",x"45",x"25",x"6d",x"92",x"6d",x"49",x"25",x"24",x"49",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"20",x"24",x"00",x"20",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"45",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6e",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"8e",x"b6"),
     (x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"96",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"49",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"24",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"45",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"db",x"92",x"69",x"6d",x"6d",x"6d",x"b6",x"49",x"6d",x"6d",x"b6",x"92",x"6d",x"6d",x"92",x"92",x"49",x"69",x"49",x"b6",x"6d",x"69",x"69",x"6d",x"b6",x"92",x"92",x"b6",x"ff",x"49",x"49",x"69",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"92",x"db",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"49",x"6d",x"b2",x"92",x"69",x"49",x"49",x"49",x"92",x"69",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"24",x"00",x"00",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"92",x"49",x"48",x"24",x"45",x"24",x"24",x"49",x"24",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"49",x"92",x"92",x"69",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"6d"),
     (x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"49",x"45",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"b6",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"92",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"25",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6e",x"8e",x"6d",x"6d",x"49",x"24",x"24",x"49",x"92",x"6d",x"24",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"69",x"92",x"92",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"6d",x"db",x"b6",x"b6",x"db",x"b6",x"69",x"6d",x"49",x"6d",x"db",x"db",x"b6",x"db",x"db",x"69",x"6d",x"6d",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"b6",x"8d",x"6d",x"92",x"ff",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6e",x"45",x"49",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"04",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"45",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"92",x"6d",x"24",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49"),
     (x"49",x"49",x"6d",x"6d",x"4d",x"92",x"db",x"ff",x"ff",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"25",x"24",x"25",x"49",x"6e",x"6e",x"49",x"24",x"45",x"49",x"45",x"24",x"49",x"49",x"49",x"b6",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"25",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"20",x"20",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"20",x"00",x"24",x"20",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"24",x"20",x"20",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"6d",x"69",x"6d",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"b6",x"db",x"69",x"6d",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"92",x"b6",x"6d",x"69",x"6d",x"6d",x"b6",x"6d",x"6d",x"92",x"b6",x"69",x"6d",x"49",x"69",x"92",x"b6",x"6d",x"69",x"6d",x"b6",x"92",x"92",x"92",x"ff",x"92",x"49",x"49",x"49",x"92",x"8e",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"25",x"25",x"25",x"25",x"6e",x"6d",x"49",x"24",x"25",x"45",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"24",x"00",x"00",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"20",x"00",x"45",x"24",x"20",x"00",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"49",x"92",x"6d",x"24",x"24",x"24",x"25",x"25",x"24",x"25",x"8e",x"92",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"25",x"24",x"24",x"25",x"25",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"db",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"25",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"49",x"45",x"24",x"24",x"49",x"49",x"92",x"b6",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"25",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"6d",x"b6",x"6d",x"69",x"69",x"6d",x"b6",x"49",x"49",x"69",x"69",x"92",x"db",x"92",x"b6",x"ff",x"6d",x"6d",x"49",x"6d",x"6d",x"db",x"b6",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"6d",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"b6",x"6d",x"49",x"6d",x"6d",x"92",x"92",x"6d",x"69",x"49",x"49",x"45",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"6d",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"00",x"24",x"69",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"25",x"49",x"b2",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"6d",x"b6",x"49",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"25",x"24",x"49",x"49",x"24",x"25",x"6d",x"92",x"6d",x"49",x"49",x"6d",x"6d",x"92",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"b6",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"6d",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"45",x"45",x"25",x"24",x"49",x"b6",x"49",x"24",x"25",x"25",x"24",x"24",x"49",x"6d",x"49",x"b6",x"92",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"49",x"45",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"25",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"25",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"20",x"00",x"49",x"49",x"24",x"24",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"49",x"45",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"fb",x"92",x"6d",x"6d",x"b6",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"69",x"6d",x"6d",x"92",x"b6",x"6d",x"6d",x"92",x"b6",x"6d",x"6d",x"6d",x"6d",x"b6",x"6d",x"6d",x"6d",x"b6",x"6d",x"69",x"6d",x"49",x"6d",x"fb",x"db",x"b2",x"b6",x"db",x"6d",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"49",x"45",x"25",x"44",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"20",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"b7",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"6d",x"49",x"49",x"24",x"45",x"24",x"24",x"49",x"db",x"6d",x"49",x"49",x"49",x"45",x"24",x"24",x"25",x"24",x"6d",x"92",x"49",x"24",x"49",x"49",x"25",x"24",x"49",x"6e",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"db",x"69",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"b2",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"25",x"49",x"49",x"49",x"25",x"49",x"b6",x"49",x"24",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"d7",x"6d",x"25",x"25",x"25",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"49",x"45",x"6d",x"92",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"6d",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"92",x"b2",x"92",x"92",x"92",x"b6",x"8e",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"6d",x"69",x"db",x"b6",x"92",x"92",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"69",x"6d",x"6d",x"69",x"d6",x"db",x"92",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6e",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"45",x"8e",x"25",x"45",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"b6",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"45",x"45",x"24",x"24",x"24",x"25",x"b6",x"92",x"48",x"49",x"49",x"45",x"44",x"24",x"24",x"24",x"69",x"b6",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"92",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"69",x"49",x"49",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b2",x"92",x"49",x"49",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"6d",x"49",x"49",x"6d",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"45",x"25",x"49",x"25",x"45",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"49",x"24",x"49",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"45",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"db",x"69",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"db",x"b6",x"b6",x"b6",x"ff",x"6d",x"49",x"69",x"69",x"69",x"b6",x"92",x"6d",x"6d",x"b6",x"92",x"49",x"69",x"6d",x"6d",x"b6",x"b6",x"92",x"92",x"ff",x"6d",x"69",x"49",x"69",x"49",x"b6",x"6d",x"49",x"49",x"49",x"92",x"db",x"92",x"92",x"92",x"b6",x"92",x"49",x"69",x"92",x"db",x"92",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"44",x"24",x"24",x"24",x"6d",x"db",x"49",x"48",x"48",x"45",x"44",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"25",x"49",x"49",x"25",x"24",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"49",x"49",x"6d",x"49",x"49",x"8e",x"b6",x"ff",x"b6",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"69",x"db",x"49",x"49",x"49",x"49"),
     (x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"4d",x"49",x"6d",x"6d",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"24",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"20",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"49",x"20",x"00",x"00",x"20",x"20",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"45",x"49",x"69",x"49",x"49",x"45",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"db",x"6d",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"d6",x"b6",x"6d",x"8e",x"b6",x"92",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"69",x"6d",x"b6",x"6d",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"69",x"49",x"6d",x"b2",x"49",x"49",x"49",x"49",x"92",x"db",x"69",x"49",x"49",x"6d",x"d7",x"b6",x"6d",x"49",x"49",x"69",x"b6",x"b6",x"49",x"49",x"49",x"49",x"92",x"92",x"25",x"25",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"25",x"69",x"db",x"6d",x"49",x"48",x"49",x"24",x"45",x"24",x"24",x"45",x"b6",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"69",x"49",x"49",x"49",x"49",x"6e",x"b6",x"db",x"fb",x"8d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"49",x"49",x"49"),
     (x"bb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"69",x"49",x"49",x"6d",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b6",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"6e",x"49",x"49",x"49",x"6d",x"6e",x"92",x"6d",x"25",x"29",x"49",x"49",x"45",x"45",x"49",x"49",x"92",x"6d",x"25",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"45",x"49",x"25",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"45",x"45",x"45",x"49",x"24",x"24",x"49",x"24",x"24",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"20",x"20",x"24",x"00",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"20",x"20",x"24",x"00",x"24",x"00",x"00",x"20",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"00",x"00",x"00",x"24",x"45",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"45",x"24",x"00",x"20",x"49",x"00",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"49",x"6e",x"92",x"25",x"49",x"49",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"92",x"b6",x"b2",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"b2",x"db",x"6d",x"69",x"6d",x"49",x"49",x"b6",x"b6",x"6d",x"92",x"b6",x"92",x"49",x"69",x"49",x"6d",x"6d",x"ff",x"b6",x"6d",x"92",x"b6",x"92",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"92",x"69",x"49",x"49",x"49",x"49",x"92",x"69",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"4d",x"49",x"24",x"24",x"24",x"49",x"49",x"b6",x"92",x"49",x"24",x"45",x"49",x"44",x"45",x"45",x"24",x"92",x"6d",x"48",x"49",x"24",x"45",x"49",x"49",x"49",x"24",x"6d",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"49",x"49",x"69",x"6d",x"b6",x"b7",x"ff",x"b6",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"d6",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"69",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"6e",x"92",x"92",x"49",x"25",x"49",x"49",x"45",x"45",x"45",x"49",x"49",x"b6",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"25",x"25",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"69",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"24",x"00",x"20",x"00",x"24",x"45",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"25",x"45",x"49",x"49",x"b6",x"6e",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"6e",x"db",x"b6",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"b6",x"b2",x"6d",x"49",x"6d",x"b6",x"6d",x"69",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"69",x"d7",x"db",x"92",x"6d",x"92",x"b6",x"6d",x"49",x"69",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"25",x"6e",x"6d",x"45",x"24",x"24",x"49",x"49",x"6d",x"69",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"00",x"00",x"24",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"45",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"25",x"49",x"49",x"6d",x"db",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"44",x"49",x"49",x"49",x"24",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"6d",x"6d",x"49",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"fb",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"6e",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"24",x"24",x"25",x"25",x"24",x"24",x"49",x"49",x"d7",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"20",x"25",x"00",x"00",x"20",x"20",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"25",x"25",x"25",x"92",x"25",x"25",x"45",x"45",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"b6",x"8e",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"db",x"b2",x"6d",x"92",x"b6",x"92",x"69",x"69",x"69",x"69",x"6d",x"ff",x"b6",x"b6",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"69",x"92",x"b6",x"92",x"8e",x"92",x"92",x"b6",x"6d",x"49",x"6d",x"6d",x"92",x"92",x"92",x"69",x"6d",x"6d",x"49",x"49",x"6d",x"b2",x"6d",x"25",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"20",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"6d",x"49",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"8e",x"6d",x"6d",x"92",x"92",x"b6",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"96",x"ff",x"d7",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"df",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"92",x"24",x"24",x"45",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"db",x"ff",x"72",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"6e",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"25",x"24",x"24",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"b6",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"25",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"24",x"24",x"24",x"45",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"b2",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"69",x"6d",x"b2",x"92",x"49",x"49",x"49",x"49",x"92",x"92",x"69",x"49",x"69",x"6d",x"b6",x"6d",x"6d",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"25",x"25",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"25",x"24",x"24",x"24",x"49",x"25",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"92",x"6e",x"92",x"92",x"92",x"92",x"b6",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"db",x"6d",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"24",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"b6",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"25",x"24",x"24",x"49",x"92",x"6d",x"24",x"25",x"49",x"45",x"49",x"49",x"49",x"44",x"92",x"92",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"25",x"24",x"24",x"00",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"20",x"24",x"6d",x"24",x"24",x"24",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6e",x"92",x"6e",x"49",x"24",x"24",x"49",x"92",x"d7",x"49",x"45",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"6d",x"92",x"92",x"6d",x"92",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"92",x"b6",x"db",x"69",x"49",x"49",x"49",x"49",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"69",x"b6",x"d7",x"6d",x"69",x"6d",x"b2",x"92",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"49",x"45",x"25",x"25",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"49",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"45",x"00",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"20",x"20",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"92",x"92",x"92",x"6d",x"6d",x"92",x"d7",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"6d",x"6d",x"49",x"69",x"49",x"49",x"69",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"db",x"ff",x"b6",x"6e",x"6d",x"49",x"49",x"6d",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"25",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8e",x"25",x"24",x"49",x"25",x"24",x"49",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"6d",x"25",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"20",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"45",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"49",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"25",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"8d",x"db",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"49",x"49",x"49",x"49",x"69",x"db",x"6d",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"6d",x"6d",x"6d",x"b6",x"6d",x"49",x"69",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"69",x"6d",x"92",x"b6",x"6d",x"6d",x"92",x"db",x"db",x"69",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"25",x"25",x"45",x"6d",x"92",x"6e",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"20",x"24",x"24",x"00",x"24",x"24",x"20",x"20",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"6d",x"49",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"20",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"44",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"b6",x"b6",x"6e",x"6d",x"49",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"6d",x"69",x"69",x"69",x"49",x"69",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"92",x"db",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b2",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6e",x"49",x"24",x"49",x"25",x"25",x"24",x"49",x"92",x"6d",x"24",x"25",x"49",x"25",x"49",x"49",x"24",x"49",x"b6",x"25",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"49",x"00",x"00",x"20",x"24",x"20",x"20",x"49",x"49",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"45",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"25",x"69",x"24",x"24",x"24",x"25",x"25",x"45",x"92",x"25",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"b6",x"b6",x"92",x"6d",x"b6",x"ff",x"6d",x"69",x"49",x"49",x"49",x"69",x"db",x"92",x"6d",x"8e",x"b6",x"92",x"49",x"69",x"49",x"49",x"49",x"db",x"db",x"92",x"b6",x"fb",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"6d",x"49",x"49",x"49",x"92",x"db",x"b2",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"8e",x"49",x"45",x"45",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"24",x"20",x"20",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"6d",x"45",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"25",x"8e",x"92",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"4d",x"49",x"49",x"49",x"45",x"49",x"45",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"8e",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"69",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"44"),
     (x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"69",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"db",x"db",x"92",x"92",x"6e",x"6e",x"6e",x"92",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"45",x"49",x"25",x"25",x"24",x"49",x"b6",x"6d",x"24",x"25",x"49",x"25",x"49",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"00",x"00",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"24",x"20",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"49",x"45",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"b2",x"b6",x"92",x"92",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"8e",x"b6",x"6d",x"6d",x"6d",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"d7",x"6d",x"49",x"49",x"69",x"92",x"b6",x"6d",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"25",x"24",x"45",x"24",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"20",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"20",x"00",x"00",x"49",x"20",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"25",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"49",x"25",x"25",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"8e",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"6d",x"db",x"db",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"44"),
     (x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"45",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"8d",x"b6",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"db",x"92",x"6d",x"6d",x"6e",x"92",x"b6",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"25",x"24",x"45",x"25",x"25",x"25",x"24",x"49",x"92",x"6d",x"24",x"25",x"49",x"49",x"25",x"24",x"49",x"92",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"49",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"69",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"92",x"92",x"49",x"45",x"45",x"49",x"92",x"b6",x"92",x"6d",x"49",x"49",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"69",x"fb",x"db",x"92",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"69",x"6d",x"92",x"92",x"49",x"49",x"6d",x"b6",x"fb",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"49",x"25",x"24",x"25",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"69",x"49",x"20",x"20",x"24",x"00",x"20",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"20",x"49",x"49",x"20",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"25",x"25",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"d6",x"ff",x"92",x"69",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24"),
     (x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"45",x"44",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"b6",x"8d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"b6",x"db",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"df",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"25",x"25",x"49",x"49",x"24",x"49",x"b6",x"6d",x"24",x"24",x"49",x"49",x"24",x"24",x"6d",x"45",x"24",x"49",x"45",x"24",x"25",x"24",x"69",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"20",x"00",x"24",x"24",x"49",x"24",x"00",x"24",x"00",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"04",x"00",x"20",x"20",x"24",x"6d",x"49",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"49",x"45",x"24",x"6d",x"92",x"45",x"49",x"45",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"db",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"b6",x"92",x"69",x"69",x"6d",x"6e",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"69",x"6d",x"92",x"b2",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"6d",x"49",x"6d",x"b6",x"8e",x"6d",x"6d",x"92",x"db",x"b6",x"69",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"45",x"45",x"49",x"6d",x"b2",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"24",x"25",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45"),
     (x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"44",x"44",x"24",x"44",x"45",x"49",x"49",x"49",x"49",x"49",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"4d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"db",x"6e",x"49",x"49",x"49",x"6d",x"92",x"db",x"db",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"24",x"25",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"20",x"20",x"45",x"24",x"00",x"20",x"00",x"00",x"24",x"20",x"00",x"00",x"20",x"24",x"20",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"45",x"25",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"92",x"b2",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"6d",x"49",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"92",x"b6",x"ff",x"8e",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"db",x"92",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"49",x"49",x"49",x"92",x"b2",x"8e",x"49",x"49",x"45",x"45",x"6d",x"b6",x"69",x"24",x"25",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"20",x"20",x"00",x"24",x"24",x"20",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"4d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92",x"d7",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"b6",x"d7",x"92",x"92",x"92",x"b6",x"b7",x"b6",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"fb",x"91",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49"),
     (x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"24",x"44",x"44",x"48",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"6d",x"49",x"69",x"6d",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"25",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"25",x"45",x"45",x"49",x"49",x"b2",x"49",x"45",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"69",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"d7",x"b2",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"69",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"69",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"45",x"45",x"25",x"25",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"20",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"24",x"24",x"25",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"6d",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"d7",x"b6",x"b2",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"69",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92"),
     (x"6d",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"45",x"24",x"44",x"44",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"6d",x"6d",x"69",x"6d",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"72",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"25",x"24",x"25",x"49",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"49",x"49",x"25",x"25",x"25",x"49",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"20",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"20",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"25",x"24",x"24",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"45",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"45",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"45",x"49",x"6d",x"92",x"92",x"92",x"6d",x"49",x"49",x"92",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"69",x"49",x"69",x"92",x"d7",x"49",x"49",x"49",x"49",x"49",x"69",x"fb",x"d7",x"8e",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"8e",x"6d",x"49",x"49",x"49",x"49",x"45",x"69",x"6d",x"25",x"25",x"24",x"24",x"25",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"6d",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"49",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"29",x"49",x"6d",x"49",x"29",x"25",x"29",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"fb",x"db",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"8d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db"),
     (x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"24",x"49",x"45",x"48",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"69",x"6d",x"6d",x"6e",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"25",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"24",x"24",x"25",x"24",x"25",x"24",x"45",x"25",x"92",x"92",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"25",x"49",x"24",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"b2",x"24",x"24",x"24",x"25",x"25",x"49",x"b6",x"6d",x"45",x"45",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"6d",x"b6",x"8e",x"69",x"69",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"b6",x"8e",x"92",x"b6",x"d7",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"6d",x"6d",x"92",x"92",x"49",x"49",x"6d",x"92",x"b6",x"b2",x"49",x"45",x"49",x"49",x"6d",x"b6",x"92",x"49",x"25",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"49",x"24",x"24",x"24",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"fb",x"db",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"df",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"d7",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"92",x"ff",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"49",x"44",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"8e",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"25",x"24",x"6d",x"b6",x"49",x"25",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"29",x"49",x"49",x"49",x"24",x"24",x"25",x"24",x"25",x"25",x"49",x"24",x"45",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"00",x"24",x"00",x"00",x"20",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"20",x"20",x"00",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"45",x"45",x"45",x"49",x"49",x"69",x"8e",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"92",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"8e",x"6d",x"6d",x"b6",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"92",x"49",x"49",x"49",x"49",x"8e",x"b6",x"92",x"6d",x"49",x"49",x"49",x"69",x"92",x"8e",x"49",x"25",x"24",x"25",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"69",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"25",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"92",x"b6",x"49",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"fb",x"b6",x"8e",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"8e",x"b6",x"ff",x"ff",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"45",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"6d",x"24",x"49",x"25",x"24",x"25",x"24",x"6d",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"25",x"24",x"24",x"24",x"49",x"72",x"29",x"24",x"25",x"24",x"24",x"49",x"45",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"44",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"20",x"20",x"24",x"24",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"00",x"20",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"24",x"25",x"49",x"45",x"49",x"45",x"b6",x"69",x"45",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"6d",x"6e",x"b6",x"92",x"49",x"49",x"49",x"49",x"69",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"b6",x"92",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"69",x"69",x"92",x"b6",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"49",x"49",x"45",x"45",x"45",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"25",x"69",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"20",x"20",x"00",x"00",x"24",x"49",x"20",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"6d",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"25",x"25",x"49",x"49",x"92",x"b7",x"49",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"6d",x"92",x"49",x"25",x"24",x"24",x"25",x"24",x"49",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"6d",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"b6",x"8d",x"6d",x"6d",x"6d",x"6e",x"b6",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"8e",x"b6",x"ff",x"ff",x"ff",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"d7",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"69"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"24",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"6d",x"6d",x"92",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"25",x"49",x"24",x"25",x"25",x"49",x"49",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"6d",x"24",x"24",x"24",x"49",x"49",x"24",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"00",x"24",x"20",x"20",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"45",x"24",x"45",x"6d",x"8e",x"92",x"6d",x"49",x"45",x"25",x"6d",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"b2",x"6d",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"d7",x"92",x"92",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"8e",x"49",x"49",x"25",x"25",x"45",x"45",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"69",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"49",x"69",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"69",x"b6",x"49",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"92",x"92",x"25",x"25",x"49",x"25",x"25",x"45",x"25",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"ff",x"b6",x"6d",x"69",x"69",x"6d",x"6d",x"72",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"ff",x"b6",x"b6",x"92",x"92",x"92",x"92",x"b7",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"69",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"25",x"24",x"45",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"45",x"49",x"24",x"00",x"20",x"24",x"25",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"b2",x"49",x"25",x"25",x"24",x"45",x"49",x"b6",x"8e",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b2",x"92",x"92",x"d7",x"fb",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"d7",x"92",x"92",x"db",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"b6",x"8e",x"92",x"8e",x"92",x"92",x"69",x"45",x"49",x"49",x"8e",x"b6",x"92",x"49",x"24",x"25",x"45",x"49",x"6d",x"92",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"45",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"45",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"49",x"45",x"20",x"24",x"24",x"20",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"6d",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"25",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"6e",x"6d",x"49",x"49",x"45",x"25",x"25",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b7",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"92",x"ff",x"b6",x"92",x"6d",x"6d",x"6e",x"b6",x"db",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"d7",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"ff",x"db",x"92",x"92",x"92",x"92",x"b2",x"b6",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"49",x"49",x"92",x"6d",x"24",x"24",x"25",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"20",x"00",x"24",x"6d",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"45",x"24",x"45",x"45",x"24",x"6d",x"6d",x"45",x"45",x"45",x"49",x"45",x"49",x"8e",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"69",x"6d",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"6d",x"b6",x"69",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"8e",x"49",x"49",x"49",x"49",x"6d",x"92",x"8e",x"6d",x"49",x"45",x"45",x"49",x"6d",x"92",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"24",x"00",x"00",x"00",x"00",x"00",x"25",x"25",x"00",x"00",x"00",x"25",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"20",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"20",x"00",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"20",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"6d",x"92",x"49",x"49",x"45",x"25",x"25",x"24",x"25",x"24",x"6d",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"db",x"db",x"92",x"8d",x"6e",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"b6",x"6d",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"69",x"69",x"69",x"6d",x"6d",x"6d",x"db",x"db",x"92",x"6e",x"92",x"92",x"b6",x"b7",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"49",x"49",x"25",x"45",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"45",x"92",x"92",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"20",x"00",x"00",x"20",x"24",x"49",x"49",x"24",x"00",x"20",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"20",x"24",x"49",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"49",x"49",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"25",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"25",x"25",x"25",x"92",x"49",x"24",x"45",x"45",x"45",x"45",x"6d",x"db",x"8e",x"49",x"49",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"8e",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"6d",x"6e",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"d7",x"92",x"92",x"b2",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"8e",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"6d",x"45",x"49",x"49",x"49",x"45",x"45",x"92",x"6d",x"45",x"25",x"24",x"24",x"24",x"45",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"49",x"49",x"45",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"6d",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"49",x"92",x"6e",x"6d",x"49",x"4d",x"6d",x"6e",x"b6",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d",x"db",x"db",x"6d",x"49",x"49",x"69",x"69",x"6d",x"6d",x"92",x"ff",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"db",x"ff",x"fb",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b7",x"ff",x"fb",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"fb",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b7",x"6d",x"69",x"49",x"6d",x"6d",x"6e",x"6d",x"45",x"24",x"45",x"25",x"45",x"45",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"4d",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"6d",x"49",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"49",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"69",x"25",x"24",x"24",x"49",x"6d",x"92",x"92",x"6d",x"49",x"45",x"49",x"92",x"6d",x"49",x"49",x"49",x"6d",x"b6",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"b2",x"6d",x"6d",x"6d",x"b2",x"db",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"b2",x"49",x"45",x"45",x"25",x"25",x"25",x"49",x"92",x"45",x"45",x"25",x"24",x"25",x"24",x"25",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"45",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"00",x"00",x"20",x"20",x"00",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"00",x"20",x"20",x"00",x"20",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"00",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"24",x"29",x"24",x"24",x"25",x"6d",x"92",x"92",x"6d",x"6d",x"49",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"69",x"6d",x"49",x"6d",x"b7",x"db",x"b6",x"92",x"b6",x"b6",x"db",x"db",x"db",x"db",x"ff",x"b6",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49"),
     (x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6e",x"6d",x"49",x"6d",x"6e",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"6d",x"6e",x"92",x"49",x"24",x"25",x"25",x"25",x"25",x"24",x"49",x"49",x"49",x"b6",x"db",x"49",x"29",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"6d",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"20",x"49",x"6d",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"20",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"25",x"24",x"20",x"24",x"24",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"25",x"49",x"69",x"92",x"8e",x"49",x"45",x"45",x"45",x"49",x"6d",x"b6",x"49",x"44",x"45",x"45",x"45",x"49",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"8e",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"6d",x"b2",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"69",x"49",x"49",x"8e",x"b2",x"b6",x"6d",x"45",x"25",x"25",x"24",x"49",x"92",x"b2",x"49",x"24",x"24",x"25",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"20",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"25",x"24",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"25",x"25",x"25",x"24",x"24",x"49",x"92",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"b6",x"b6",x"b6",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"6d",x"69",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"d7",x"6d",x"49",x"49",x"49",x"49"),
     (x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"d7",x"b6",x"4d",x"49",x"49",x"49",x"6d",x"b6",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"b6",x"b7",x"4d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"25",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"49",x"b6",x"b6",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"24",x"49",x"24",x"24",x"49",x"49",x"45",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"00",x"00",x"00",x"24",x"24",x"00",x"24",x"20",x"00",x"20",x"24",x"20",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"25",x"45",x"45",x"45",x"45",x"6d",x"6d",x"45",x"45",x"45",x"49",x"49",x"49",x"69",x"b2",x"49",x"45",x"45",x"45",x"49",x"8e",x"92",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"b2",x"8e",x"6d",x"6d",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"8e",x"8e",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"45",x"25",x"49",x"6d",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"45",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"20",x"00",x"00",x"20",x"24",x"6d",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"25",x"25",x"24",x"25",x"6d",x"db",x"49",x"49",x"49",x"49",x"45",x"45",x"25",x"25",x"24",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"ff",x"db",x"db",x"db",x"d7",x"b6",x"92",x"92",x"db",x"db",x"b6",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"92",x"49",x"49",x"25",x"25",x"49",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"49",x"25",x"49",x"45",x"45",x"49",x"49",x"92",x"92",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"24",x"49",x"45",x"24",x"24",x"49",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"45",x"24",x"24",x"24",x"25",x"49",x"00",x"00",x"00",x"20",x"20",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"6d",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"25",x"25",x"24",x"45",x"92",x"49",x"45",x"45",x"45",x"45",x"45",x"92",x"b6",x"92",x"8e",x"6e",x"92",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"8e",x"49",x"49",x"6d",x"b2",x"d7",x"49",x"49",x"49",x"45",x"45",x"45",x"49",x"92",x"69",x"45",x"45",x"45",x"45",x"45",x"45",x"6d",x"92",x"49",x"25",x"45",x"25",x"25",x"25",x"69",x"b2",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"25",x"24",x"24",x"24",x"25",x"25",x"20",x"00",x"20",x"20",x"20",x"00",x"20",x"24",x"25",x"24",x"20",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"45",x"24",x"24",x"00",x"00",x"00",x"00",x"20",x"49",x"6d",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"b6",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"4d",x"49",x"25",x"24",x"24",x"24",x"45",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"d6",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"df",x"71",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"45",x"49",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"69",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"b2",x"49",x"24",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"24",x"24",x"25",x"25",x"45",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"44",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"20",x"00",x"24",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"25",x"6d",x"92",x"8e",x"8e",x"6d",x"6d",x"8e",x"b2",x"49",x"49",x"45",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"d7",x"b6",x"92",x"92",x"92",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"8e",x"49",x"49",x"69",x"8e",x"92",x"49",x"45",x"45",x"49",x"49",x"8e",x"b2",x"45",x"49",x"45",x"45",x"45",x"45",x"25",x"92",x"49",x"25",x"25",x"24",x"25",x"25",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"49",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"25",x"6d",x"25",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"6e",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"8e",x"b6",x"49",x"44",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"25",x"49",x"49",x"6d",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"6e",x"92",x"db",x"db",x"b6",x"92",x"8e",x"6d",x"6d",x"6d",x"6e",x"db",x"ff",x"ff",x"fb",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6e",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"69",x"92",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"25",x"49",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"25",x"24",x"25",x"49",x"92",x"6d",x"24",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"b2",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"25",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"25",x"45",x"25",x"25",x"49",x"92",x"8e",x"45",x"25",x"45",x"45",x"45",x"49",x"49",x"92",x"6d",x"45",x"45",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"69",x"45",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"b6",x"92",x"8e",x"6d",x"8e",x"92",x"6d",x"49",x"45",x"45",x"45",x"49",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"25",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"45",x"49",x"20",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"00",x"00",x"24",x"49",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"49",x"49",x"24",x"24",x"24",x"00",x"24",x"00",x"00",x"25",x"6d",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"25",x"49",x"6e",x"b6",x"49",x"49",x"45",x"49",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"25",x"92",x"96",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6e",x"b6",x"db",x"d7",x"92",x"92",x"8e",x"6e",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"69",x"6d",x"b6",x"ff",x"ff",x"b7",x"8e",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"25",x"24",x"24",x"49",x"92",x"6d",x"24",x"25",x"45",x"49",x"49",x"24",x"24",x"49",x"6d",x"92",x"25",x"24",x"49",x"49",x"25",x"45",x"25",x"92",x"92",x"45",x"24",x"24",x"25",x"45",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"00",x"20",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"00",x"24",x"49",x"25",x"24",x"20",x"24",x"24",x"25",x"49",x"00",x"00",x"20",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"25",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"45",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"49",x"24",x"24",x"24",x"25",x"24",x"25",x"45",x"92",x"49",x"24",x"25",x"45",x"45",x"45",x"49",x"92",x"b6",x"92",x"8e",x"6d",x"92",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"6d",x"6d",x"6d",x"b2",x"d7",x"69",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"45",x"49",x"45",x"45",x"49",x"b2",x"92",x"8e",x"6d",x"49",x"49",x"6d",x"8e",x"69",x"45",x"45",x"49",x"6d",x"6d",x"6e",x"92",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"45",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"25",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"49",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"6e",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"25",x"49",x"6d",x"d7",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"92",x"8e",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6e",x"92",x"b6",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"24",x"49",x"25",x"24",x"49",x"92",x"b2",x"49",x"25",x"49",x"49",x"49",x"24",x"49",x"49",x"6d",x"6d",x"24",x"25",x"49",x"45",x"24",x"25",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"20",x"24",x"00",x"24",x"00",x"00",x"00",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"20",x"24",x"24",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"6d",x"b6",x"6d",x"49",x"45",x"25",x"49",x"8e",x"6d",x"45",x"49",x"49",x"49",x"49",x"8e",x"8e",x"45",x"49",x"49",x"45",x"45",x"49",x"49",x"b2",x"6d",x"49",x"49",x"49",x"49",x"8e",x"92",x"49",x"45",x"45",x"45",x"45",x"49",x"92",x"6d",x"45",x"45",x"25",x"25",x"25",x"25",x"45",x"92",x"6d",x"45",x"45",x"45",x"45",x"45",x"24",x"6d",x"b6",x"6e",x"49",x"24",x"24",x"24",x"25",x"49",x"6e",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"25",x"6d",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"00",x"00",x"24",x"20",x"00",x"20",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"24",x"24",x"25",x"49",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"25",x"24",x"25",x"49",x"6e",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"6e",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"6d",x"92",x"ff",x"ff",x"b6",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"db",x"6d",x"49",x"49",x"49",x"69",x"6d",x"69",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"b6",x"92",x"6e",x"8e",x"92",x"b6",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"49",x"25",x"49",x"49",x"92",x"49",x"25",x"49",x"25",x"24",x"49",x"6d",x"49",x"6d",x"49",x"24",x"49",x"49",x"49",x"24",x"49",x"49",x"49",x"b7",x"6d",x"25",x"24",x"24",x"25",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"25",x"92",x"49",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"45",x"92",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"20",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"25",x"6d",x"8e",x"69",x"49",x"49",x"6d",x"8e",x"b6",x"6d",x"45",x"45",x"45",x"45",x"49",x"49",x"49",x"8e",x"6e",x"49",x"45",x"45",x"45",x"49",x"92",x"49",x"45",x"45",x"49",x"45",x"45",x"45",x"49",x"b6",x"92",x"6d",x"6d",x"92",x"b6",x"b6",x"49",x"45",x"45",x"45",x"25",x"25",x"25",x"49",x"92",x"25",x"45",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"00",x"00",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"6d",x"49",x"24",x"24",x"49",x"b6",x"6d",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"25",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"92",x"b6",x"49",x"49",x"49",x"29",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"b7",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"8e",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"db",x"b6",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"d6",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"24",x"24",x"25",x"25",x"49",x"49",x"49",x"b6",x"6d",x"25",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"24",x"45",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"b6",x"6d",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"25",x"04",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"20",x"20",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6e",x"b2",x"49",x"24",x"24",x"25",x"24",x"24",x"45",x"69",x"92",x"45",x"25",x"25",x"45",x"25",x"25",x"45",x"6d",x"b6",x"92",x"6e",x"6d",x"92",x"b6",x"92",x"45",x"49",x"49",x"45",x"45",x"25",x"45",x"49",x"b2",x"6d",x"49",x"45",x"45",x"49",x"49",x"8e",x"6d",x"45",x"45",x"45",x"49",x"6d",x"b6",x"6d",x"25",x"24",x"24",x"24",x"49",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"20",x"24",x"25",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"25",x"49",x"49",x"24",x"24",x"24",x"8e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"25",x"25",x"92",x"92",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"6d",x"92",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"fb",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"db",x"92",x"6d",x"69",x"6d",x"6d",x"92",x"b6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"6e",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"25",x"49",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"b6",x"6e",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"00",x"24",x"24",x"20",x"00",x"49",x"69",x"49",x"24",x"24",x"25",x"49",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"69",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"92",x"49",x"25",x"24",x"24",x"25",x"24",x"24",x"45",x"6d",x"8e",x"45",x"25",x"25",x"25",x"45",x"6d",x"8e",x"49",x"45",x"45",x"25",x"45",x"49",x"6d",x"6d",x"45",x"25",x"45",x"25",x"24",x"45",x"92",x"69",x"45",x"45",x"45",x"25",x"45",x"45",x"49",x"92",x"b6",x"6e",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"45",x"6d",x"92",x"b2",x"6d",x"24",x"24",x"25",x"24",x"24",x"49",x"8e",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"20",x"20",x"25",x"24",x"20",x"00",x"00",x"00",x"20",x"49",x"49",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"20",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"24",x"20",x"00",x"00",x"24",x"24",x"20",x"00",x"00",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"49",x"25",x"49",x"49",x"45",x"24",x"24",x"49",x"6e",x"25",x"24",x"24",x"49",x"45",x"25",x"45",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"6e",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"b7",x"db",x"b6",x"b6",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"49",x"49",x"69",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"8e",x"49",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"b6",x"6e",x"6d",x"6d",x"6e",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"6e",x"49",x"45",x"49",x"49",x"49",x"49",x"8e",x"6d",x"25",x"25",x"49",x"49",x"49",x"25",x"25",x"24",x"49",x"b6",x"92",x"49",x"25",x"25",x"45",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"20",x"24",x"00",x"24",x"45",x"24",x"00",x"20",x"00",x"00",x"00",x"20",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"92",x"6d",x"6d",x"8e",x"b2",x"b2",x"49",x"45",x"45",x"45",x"45",x"45",x"25",x"45",x"8e",x"b2",x"6d",x"6d",x"6d",x"8e",x"b6",x"92",x"45",x"45",x"49",x"45",x"25",x"45",x"24",x"45",x"92",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"25",x"45",x"45",x"49",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"45",x"25",x"49",x"69",x"6e",x"6e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"00",x"24",x"24",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"00",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"20",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"6d",x"49",x"25",x"25",x"49",x"49",x"45",x"25",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"25",x"24",x"24",x"25",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"45",x"45",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"b6",x"92",x"92",x"6e",x"6e",x"92",x"92",x"db",x"b6",x"6d",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b2",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"ff",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"6d"),
     (x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"db",x"6d",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"b7",x"92",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"b7",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"92",x"49",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"45",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"49",x"20",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"20",x"49",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"45",x"25",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"8e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"69",x"49",x"24",x"25",x"49",x"8e",x"69",x"25",x"25",x"25",x"25",x"25",x"49",x"92",x"49",x"45",x"24",x"24",x"25",x"24",x"45",x"45",x"8e",x"6d",x"49",x"49",x"45",x"45",x"49",x"8e",x"6d",x"45",x"24",x"25",x"24",x"24",x"45",x"6e",x"6d",x"25",x"24",x"24",x"24",x"24",x"25",x"45",x"45",x"92",x"49",x"25",x"24",x"25",x"24",x"24",x"24",x"45",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"49",x"25",x"24",x"00",x"24",x"24",x"24",x"20",x"24",x"20",x"20",x"00",x"00",x"00",x"6d",x"6d",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"6d",x"49",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"b7",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"24",x"24",x"49",x"49",x"25",x"24",x"25",x"49",x"25",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"8e",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6e",x"b6",x"db",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6"),
     (x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"71",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"da",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"db",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"6d",x"db",x"b7",x"6d",x"49",x"49",x"6d",x"92",x"b6",x"b7",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"24",x"25",x"49",x"49",x"25",x"24",x"25",x"24",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"24",x"29",x"25",x"49",x"69",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"92",x"69",x"45",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"25",x"49",x"49",x"6d",x"b6",x"6d",x"24",x"45",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"69",x"45",x"24",x"25",x"24",x"49",x"8e",x"49",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"8e",x"6d",x"6d",x"6d",x"92",x"b6",x"6d",x"25",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"45",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"20",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"49",x"44",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"24",x"24",x"45",x"b6",x"92",x"49",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"25",x"6e",x"6d",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"6d",x"92",x"b6",x"8e",x"69",x"49",x"49",x"6d",x"92",x"fb",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"6d",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"db",x"d7",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"db",x"ff",x"da",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"fb",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db"),
     (x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"db",x"b6",x"6e",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"92",x"d7",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"29",x"24",x"24",x"49",x"45",x"25",x"45",x"25",x"49",x"49",x"b6",x"b6",x"49",x"25",x"25",x"24",x"25",x"49",x"92",x"6d",x"24",x"45",x"45",x"49",x"49",x"49",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"25",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"00",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"25",x"49",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"25",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"45",x"25",x"49",x"6d",x"49",x"25",x"24",x"24",x"49",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"25",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"8e",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"25",x"24",x"25",x"24",x"25",x"24",x"25",x"24",x"49",x"92",x"69",x"45",x"25",x"24",x"24",x"45",x"6d",x"6e",x"49",x"24",x"24",x"49",x"49",x"92",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"69",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"00",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"48",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"25",x"24",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"db",x"db",x"db",x"db",x"db",x"b7",x"b7",x"db",x"ff",x"da",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"db",x"ff",x"fb",x"92",x"6d",x"6d",x"6d",x"49",x"69",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"92"),
     (x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"6d",x"92",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"49",x"45",x"49",x"49",x"49",x"49",x"b7",x"92",x"25",x"24",x"24",x"24",x"25",x"49",x"92",x"92",x"49",x"25",x"49",x"25",x"49",x"25",x"49",x"49",x"6d",x"25",x"24",x"25",x"24",x"25",x"49",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"20",x"24",x"00",x"00",x"20",x"00",x"20",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"20",x"20",x"20",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"20",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"45",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"24",x"24",x"25",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"b6",x"92",x"6d",x"49",x"49",x"45",x"49",x"6d",x"6d",x"49",x"25",x"45",x"49",x"69",x"6d",x"8e",x"8e",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"20",x"24",x"00",x"24",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"49",x"45",x"45",x"49",x"49",x"25",x"24",x"49",x"49",x"49",x"25",x"25",x"25",x"45",x"49",x"d7",x"92",x"49",x"49",x"49",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"69",x"49",x"49",x"49",x"49",x"69",x"49",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"b7",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"b6",x"b7",x"db",x"fb",x"92",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b2",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"fb",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"6d",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"24",x"24",x"49",x"25",x"25",x"49",x"49",x"92",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"6d",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"04",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"25",x"49",x"25",x"25",x"45",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6e",x"6d",x"6d",x"6d",x"8e",x"b2",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"69",x"92",x"6d",x"49",x"49",x"6d",x"8e",x"b2",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"24",x"24",x"45",x"24",x"45",x"6d",x"6e",x"8e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"25",x"24",x"25",x"49",x"25",x"24",x"20",x"20",x"20",x"20",x"20",x"20",x"20",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"8e",x"6d",x"24",x"25",x"49",x"49",x"24",x"45",x"49",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"92",x"49",x"45",x"25",x"24",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"49",x"6e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"d6",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"db",x"fb",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"28",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"91",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"91",x"b6",x"db",x"92",x"6d",x"6d",x"49",x"49",x"49",x"92",x"db",x"ff",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"25",x"24",x"25",x"49",x"6e",x"92",x"49",x"25",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"25",x"49",x"24",x"45",x"45",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"20",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"20",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"6d",x"8e",x"49",x"45",x"25",x"25",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"20",x"20",x"24",x"00",x"20",x"20",x"24",x"49",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"20",x"20",x"20",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"49",x"49",x"24",x"45",x"49",x"49",x"25",x"25",x"6d",x"6d",x"49",x"25",x"25",x"25",x"49",x"49",x"b6",x"92",x"49",x"45",x"45",x"24",x"45",x"45",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"69",x"49",x"69",x"69",x"6d",x"49",x"8e",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"92",x"49",x"49"),
     (x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"b6",x"db",x"49",x"28",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"da",x"d6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"45",x"49",x"24",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"6d",x"25",x"24",x"25",x"45",x"49",x"49",x"49",x"25",x"24",x"45",x"49",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"49",x"49",x"20",x"00",x"24",x"49",x"24",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"00",x"20",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"8e",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"49",x"45",x"49",x"49",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"8e",x"49",x"49",x"49",x"6d",x"8e",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"20",x"20",x"20",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"20",x"00",x"00",x"20",x"24",x"20",x"24",x"24",x"00",x"00",x"49",x"6d",x"49",x"24",x"24",x"20",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"25",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"24",x"49",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"92",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"49",x"6e",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"6d",x"49",x"6d",x"6d",x"6d",x"69",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"ff",x"b6",x"92",x"8d",x"8d",x"8d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"8d",x"ff",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49"),
     (x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"da",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"6d",x"25",x"45",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"25",x"49",x"49",x"24",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"20",x"00",x"00",x"00",x"24",x"20",x"20",x"20",x"24",x"24",x"00",x"20",x"00",x"00",x"00",x"20",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"49",x"69",x"6e",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"69",x"49",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"20",x"00",x"00",x"00",x"24",x"25",x"24",x"00",x"00",x"00",x"20",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"00",x"24",x"49",x"49",x"24",x"20",x"24",x"20",x"24",x"24",x"00",x"00",x"20",x"25",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"24",x"49",x"25",x"24",x"25",x"8d",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"92",x"b6",x"49",x"24",x"24",x"25",x"24",x"25",x"24",x"24",x"24",x"49",x"92",x"6e",x"49",x"49",x"25",x"25",x"49",x"49",x"b6",x"b6",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"69",x"69",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"6e",x"72",x"92",x"b6",x"ff",x"b6",x"92",x"92",x"8d",x"91",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49"),
     (x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"db",x"ff",x"fb",x"92",x"6d",x"6d",x"6d",x"6d",x"8d",x"92",x"b6",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"db",x"b6",x"49",x"25",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"00",x"24",x"20",x"20",x"00",x"00",x"00",x"24",x"20",x"24",x"25",x"25",x"24",x"24",x"24",x"45",x"69",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"92",x"92",x"8e",x"6d",x"49",x"49",x"45",x"49",x"49",x"69",x"49",x"25",x"24",x"49",x"49",x"6d",x"6d",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"45",x"49",x"49",x"69",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"25",x"49",x"49",x"24",x"00",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"25",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"44",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"49",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"69",x"b6",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"25",x"24",x"25",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"db",x"b6",x"6e",x"6d",x"6d",x"6e",x"92",x"db",x"db",x"92",x"92",x"8d",x"92",x"6d",x"6d",x"92",x"d7",x"ff",x"ff",x"db",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"92",x"49",x"49",x"49",x"49"),
     (x"db",x"92",x"6d",x"49",x"49",x"49",x"69",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"4d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"db",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"b6",x"72",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"29",x"25",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"b6",x"b6",x"49",x"24",x"24",x"24",x"45",x"24",x"49",x"92",x"92",x"49",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"24",x"49",x"24",x"24",x"00",x"00",x"20",x"24",x"25",x"25",x"20",x"20",x"24",x"24",x"24",x"20",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"6d",x"49",x"49",x"49",x"6d",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"45",x"24",x"25",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"00",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"25",x"25",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"92",x"49",x"49",x"49",x"25",x"25",x"25",x"49",x"49",x"24",x"6d",x"b6",x"6d",x"24",x"25",x"49",x"45",x"25",x"25",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"ff",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"ff",x"b6",x"92",x"92",x"92",x"8d",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49"),
     (x"ff",x"db",x"92",x"6d",x"6d",x"49",x"69",x"69",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"6d",x"b6",x"ff",x"ff",x"db",x"b6",x"8d",x"6d",x"6d",x"8d",x"92",x"da",x"db",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"92",x"92",x"25",x"24",x"24",x"45",x"49",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"45",x"69",x"8e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6e",x"69",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"20",x"24",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"49",x"24",x"20",x"00",x"00",x"24",x"49",x"6d",x"49",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"6d",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"25",x"6d",x"6d",x"24",x"49",x"45",x"45",x"49",x"49",x"49",x"25",x"92",x"92",x"49",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6e",x"92",x"ff",x"db",x"b2",x"92",x"92",x"92",x"6d",x"92",x"b6",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"8d",x"fb",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"d6",x"ff",x"ff",x"db",x"b6",x"92",x"8d",x"6d",x"92",x"b6",x"db",x"db",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"25",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"25",x"6e",x"b6",x"49",x"49",x"25",x"25",x"24",x"24",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"49",x"24",x"00",x"24",x"20",x"24",x"24",x"20",x"24",x"20",x"20",x"45",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"45",x"49",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"20",x"20",x"24",x"20",x"00",x"00",x"00",x"20",x"49",x"49",x"24",x"20",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"25",x"24",x"49",x"8e",x"49",x"24",x"25",x"25",x"49",x"25",x"25",x"49",x"92",x"6d",x"49",x"25",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"db",x"92",x"92",x"92",x"b2",x"db",x"ff",x"ff",x"db",x"6d",x"6d",x"6d",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"92",x"8d",x"92",x"b6",x"ff",x"ff",x"ff",x"db",x"91",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"db",x"fb",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"91",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"91",x"db",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"b6",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"69",x"db",x"92",x"28",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"49",x"92",x"49",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"49",x"49",x"25",x"24",x"24",x"45",x"49",x"49",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6e",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"49",x"45",x"49",x"6d",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6e",x"69",x"49",x"49",x"45",x"45",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"20",x"24",x"20",x"24",x"24",x"20",x"24",x"45",x"49",x"24",x"00",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"69",x"49",x"45",x"24",x"24",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"25",x"24",x"49",x"8e",x"49",x"24",x"25",x"24",x"25",x"25",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"25",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"b2",x"b6",x"92",x"b6",x"db",x"ff",x"ff",x"92",x"6d",x"6d",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"b6",x"ff",x"b6",x"b2",x"92",x"92",x"8e",x"92",x"b6",x"ff",x"ff",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"b6",x"ff",x"b2",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"db",x"db",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"4d",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"25",x"25",x"49",x"49",x"49",x"45",x"45",x"49",x"49",x"92",x"25",x"24",x"49",x"49",x"45",x"49",x"49",x"45",x"25",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"8e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"20",x"00",x"24",x"24",x"24",x"00",x"20",x"20",x"20",x"24",x"49",x"24",x"20",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"45",x"25",x"45",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"20",x"20",x"24",x"24",x"20",x"24",x"00",x"24",x"25",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"6d",x"6d",x"45",x"24",x"24",x"20",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"6d",x"49",x"92",x"49",x"49",x"44",x"24",x"24",x"45",x"24",x"49",x"6d",x"69",x"49",x"45",x"24",x"25",x"25",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"25",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"92",x"6d",x"6d",x"69",x"6d",x"6d",x"49",x"49",x"49",x"49",x"8e",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"b6",x"8d",x"8d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"b2",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"92",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b7",x"92",x"92",x"92",x"92",x"db",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"92",x"6d",x"49",x"49",x"49",x"6d",x"92",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"25",x"25",x"29",x"49",x"92",x"6d",x"25",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"24",x"24",x"49",x"45",x"45",x"45",x"45",x"24",x"24",x"25",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"69",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"8e",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6e",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"25",x"24",x"20",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"69",x"49",x"24",x"25",x"24",x"49",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"92",x"92",x"49",x"49",x"45",x"25",x"25",x"24",x"49",x"6d",x"6d",x"49",x"49",x"25",x"25",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"49",x"25",x"29",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"db",x"92",x"8e",x"6d",x"6d",x"92",x"b6",x"ff",x"b6",x"6d",x"6d",x"69",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"db",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"b6",x"b2",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"69",x"69",x"49",x"92",x"fb",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"49",x"49",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"b6",x"6e",x"6d",x"6d",x"92",x"db",x"db",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6e",x"6d",x"6d",x"6d",x"92",x"92",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"25",x"25",x"25",x"25",x"25",x"49",x"6d",x"92",x"49",x"49",x"45",x"49",x"49",x"49",x"45",x"45",x"49",x"69",x"24",x"24",x"25",x"45",x"49",x"49",x"25",x"25",x"25",x"49",x"6d",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"00",x"00",x"24",x"20",x"20",x"24",x"24",x"20",x"00",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"00",x"24",x"00",x"24",x"24",x"20",x"20",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"69",x"49",x"69",x"6d",x"8e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"25",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"00",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"45",x"45",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"6d",x"49",x"49",x"44",x"49",x"24",x"24",x"49",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"4d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"92",x"6d",x"69",x"6d",x"6d",x"92",x"db",x"d6",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"6d",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"fb",x"92",x"8e",x"8d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44"),
     (x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"49",x"49",x"69",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"91",x"db",x"ff",x"ff",x"db",x"db",x"db",x"b7",x"b6",x"db",x"ff",x"ff",x"92",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b7",x"92",x"6d",x"49",x"6d",x"6d",x"b6",x"db",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"b6",x"6e",x"6d",x"6d",x"6d",x"6e",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"45",x"49",x"49",x"25",x"49",x"49",x"49",x"24",x"49",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"00",x"25",x"49",x"24",x"00",x"00",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"6d",x"49",x"49",x"25",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"6d",x"92",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"b6",x"6d",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"45",x"24",x"25",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"25",x"49",x"92",x"92",x"6d",x"49",x"49",x"49",x"6d",x"6e",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"ff",x"db",x"91",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"d6",x"b2",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"6d",x"d6",x"ff",x"b2",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24"),
     (x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"6d",x"6d",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"fb",x"b6",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"25",x"25",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"25",x"24",x"25",x"25",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"8e",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"20",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"25",x"45",x"45",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"6e",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"b2",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"45",x"24",x"24",x"92",x"49",x"24",x"25",x"25",x"25",x"49",x"49",x"25",x"24",x"24",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6e",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"db",x"92",x"69",x"49",x"49",x"49",x"49",x"4d",x"92",x"db",x"92",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"8e",x"db",x"ff",x"db",x"b6",x"b6",x"b2",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"d6",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"b6",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24"),
     (x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"ff",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"6d",x"69",x"6d",x"6d",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"db",x"b6",x"b6",x"b7",x"db",x"ff",x"ff",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"6e",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6e",x"24",x"25",x"49",x"49",x"49",x"25",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"45",x"49",x"49",x"49",x"49",x"4d",x"49",x"24",x"45",x"49",x"49",x"45",x"25",x"25",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"00",x"20",x"49",x"49",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"6d",x"6d",x"49",x"49",x"6d",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"25",x"45",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"20",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"92",x"92",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b2",x"92",x"49",x"49",x"49",x"49",x"25",x"45",x"45",x"49",x"24",x"24",x"6d",x"69",x"49",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"b6",x"b6",x"49",x"49",x"25",x"24",x"25",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6e",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b2",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"db",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"92",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24"),
     (x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"6e",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"91",x"db",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"b6",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"6d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"49",x"25",x"49",x"45",x"45",x"25",x"25",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"20",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6e",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"20",x"00",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"69",x"6d",x"49",x"49",x"49",x"49",x"45",x"25",x"24",x"24",x"6d",x"92",x"49",x"49",x"44",x"49",x"24",x"24",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"49",x"92",x"92",x"6e",x"49",x"49",x"49",x"49",x"6e",x"db",x"db",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"8d",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"92",x"db",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49"),
     (x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"ff",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"6d",x"db",x"92",x"49",x"49",x"25",x"24",x"24",x"25",x"49",x"6d",x"6e",x"49",x"24",x"24",x"25",x"25",x"25",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"20",x"00",x"00",x"24",x"49",x"45",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6e",x"6d",x"49",x"49",x"45",x"45",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"00",x"00",x"24",x"24",x"20",x"24",x"24",x"00",x"00",x"00",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6e",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"49",x"25",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"49",x"49",x"49",x"49",x"24",x"25",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"24",x"24",x"25",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"24",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"fb",x"db",x"b6",x"d6",x"db",x"fb",x"ff",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"6d",x"6d",x"91",x"6d",x"6d",x"69",x"6d",x"db",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"92"),
     (x"b6",x"b6",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"24",x"44",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"db",x"92",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"fb",x"db",x"92",x"92",x"92",x"92",x"92",x"b7",x"ff",x"ff",x"ff",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"db",x"8e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d7",x"92",x"49",x"25",x"24",x"24",x"25",x"49",x"49",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"20",x"20",x"20",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"6d",x"6d",x"49",x"49",x"49",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"69",x"49",x"24",x"20",x"20",x"24",x"69",x"6d",x"69",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"49",x"49",x"24",x"24",x"49",x"6d",x"49",x"49",x"49",x"24",x"25",x"25",x"49",x"92",x"b2",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"49",x"25",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"25",x"45",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"8e",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"91",x"6d",x"6d",x"6d",x"6d",x"d7",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"24",x"92",x"92"),
     (x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"92",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"92",x"49",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"25",x"29",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"45",x"24",x"24",x"20",x"20",x"24",x"24",x"25",x"45",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"45",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"45",x"49",x"25",x"24",x"20",x"24",x"6d",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"92",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"25",x"49",x"49",x"6d",x"b7",x"92",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"49",x"24",x"6d",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"6d",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b7",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"fb",x"ff",x"db",x"92",x"92",x"6d",x"6d",x"8d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"6d",x"b6",x"6d"),
     (x"b6",x"b6",x"b6",x"b7",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8d",x"db",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"b7",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6e",x"49",x"24",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"25",x"24",x"45",x"49",x"49",x"45",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"49",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"00",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"69",x"49",x"25",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"45",x"24",x"25",x"25",x"24",x"45",x"6d",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"48",x"49",x"49",x"49",x"24",x"25",x"49",x"49",x"24",x"49",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"ff",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"ff",x"fb",x"b6",x"92",x"6d",x"6d",x"8d",x"92",x"6d",x"6d",x"6d",x"b6",x"ff",x"fb",x"8d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"6d",x"49"),
     (x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"24",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"db",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"db",x"92",x"6d",x"6d",x"69",x"49",x"6d",x"92",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"69",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"6e",x"49",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6e",x"25",x"24",x"49",x"49",x"49",x"25",x"49",x"49",x"45",x"49",x"b6",x"b6",x"49",x"25",x"24",x"24",x"24",x"25",x"24",x"24",x"49",x"8e",x"92",x"6d",x"49",x"45",x"45",x"24",x"24",x"24",x"24",x"24",x"49",x"8e",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"6d",x"24",x"00",x"00",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"20",x"24",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"25",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"69",x"49",x"49",x"49",x"69",x"6d",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"45",x"24",x"24",x"45",x"45",x"49",x"49",x"24",x"24",x"45",x"49",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"49",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"25",x"24",x"25",x"25",x"24",x"45",x"49",x"24",x"24",x"49",x"49",x"24",x"25",x"49",x"45",x"25",x"24",x"24",x"24",x"69",x"92",x"6e",x"49",x"25",x"24",x"25",x"49",x"49",x"6d",x"b6",x"b6",x"49",x"44",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"d7",x"8d",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"db",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"72",x"db",x"ff",x"ff",x"ff",x"db",x"db",x"db",x"db",x"b7",x"db",x"ff",x"ff",x"b6",x"92",x"8d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"fb",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"92",x"92",x"49",x"49"),
     (x"db",x"bb",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"fb",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"48",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"db",x"6d",x"49",x"69",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"92",x"b7",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"91",x"fb",x"b6",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"b6",x"6d",x"49",x"49",x"4d",x"6d",x"72",x"92",x"92",x"49",x"29",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"24",x"25",x"49",x"92",x"b7",x"69",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"b6",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"45",x"6d",x"49",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"49",x"49",x"49",x"24",x"24",x"49",x"25",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"25",x"25",x"25",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"49",x"6d",x"db",x"92",x"49",x"44",x"44",x"49",x"49",x"49",x"25",x"49",x"49",x"24",x"49",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"db",x"ff",x"ff",x"92",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"db",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"24",x"92",x"b6",x"49",x"49",x"45"),
     (x"ff",x"db",x"b7",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"db",x"ff",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"44",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"db",x"6d",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"fb",x"db",x"8e",x"6d",x"69",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"25",x"49",x"49",x"49",x"45",x"49",x"6d",x"6d",x"b6",x"6d",x"24",x"25",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"69",x"b6",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"b6",x"4d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6e",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"45",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"25",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"25",x"6d",x"92",x"6d",x"49",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"6d",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"49",x"49",x"24",x"49",x"6d",x"92",x"49",x"49",x"49",x"49",x"45",x"49",x"49",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"ff",x"ff",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"4d",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"91",x"6d",x"6d",x"92",x"db",x"ff",x"da",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"da",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"6d",x"b6",x"6d",x"49",x"45",x"49"),
     (x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"6d",x"24",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"b6",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"d7",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"ff",x"ff",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b2",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"b6",x"6d",x"49",x"45",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"6d",x"25",x"49",x"49",x"49",x"45",x"49",x"49",x"45",x"49",x"69",x"49",x"92",x"6d",x"24",x"25",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"92",x"6e",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"49",x"25",x"45",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"6d",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b2",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"b6",x"ff",x"db",x"b6",x"b6",x"92",x"b6",x"db",x"ff",x"ff",x"ff",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"6d",x"6d",x"92",x"ff",x"ff",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"b7",x"ff",x"db",x"b6",x"91",x"6d",x"6d",x"91",x"92",x"6d",x"6d",x"6d",x"db",x"ff",x"db",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49"),
     (x"b6",x"ff",x"ff",x"db",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"db",x"b6",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"8d",x"d7",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"92",x"6d",x"6d",x"6e",x"92",x"b7",x"ff",x"b6",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"db",x"72",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"6d",x"25",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"25",x"24",x"45",x"49",x"24",x"24",x"49",x"b6",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"49",x"6d",x"92",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"6d",x"49",x"25",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"45",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"20",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"00",x"00",x"00",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"b2",x"8e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"25",x"6d",x"6d",x"49",x"49",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"49",x"49",x"49",x"92",x"b7",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"6d",x"92",x"6d",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"6d",x"6d",x"4d",x"49",x"49",x"49",x"49",x"6d",x"d7",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"db",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"db",x"db",x"b6",x"b6",x"db",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"4d",x"4d",x"92",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"ff",x"db",x"b6",x"92",x"6d",x"6d",x"8d",x"92",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"24",x"b2",x"b2",x"49",x"49",x"45",x"49",x"49"),
     (x"b6",x"da",x"ff",x"ff",x"db",x"b7",x"b7",x"db",x"db",x"ff",x"fb",x"db",x"db",x"fb",x"ff",x"db",x"b6",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"db",x"ff",x"b6",x"6d",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"8d",x"b6",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"ff",x"92",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"b6",x"6d",x"6d",x"4d",x"6d",x"6d",x"92",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"db",x"6d",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"6d",x"49",x"24",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6e",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"69",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"6d",x"92",x"6d",x"24",x"24",x"45",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"69",x"49",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"69",x"49",x"45",x"24",x"24",x"24",x"49",x"49",x"49",x"45",x"24",x"24",x"00",x"00",x"20",x"20",x"20",x"24",x"49",x"6e",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"92",x"b6",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"25",x"25",x"6d",x"92",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"25",x"24",x"45",x"24",x"24",x"24",x"24",x"49",x"6d",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"92",x"69",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"6d",x"6e",x"6d",x"6d",x"4d",x"4d",x"6d",x"6d",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"45",x"49",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"db",x"b2",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"ff",x"db",x"db",x"db",x"b6",x"db",x"db",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"b6",x"db",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"24",x"92",x"b6",x"49",x"49",x"45",x"49",x"49",x"49"),
     (x"92",x"b6",x"db",x"ff",x"db",x"db",x"b7",x"db",x"db",x"ff",x"ff",x"db",x"db",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"df",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"ff",x"ff",x"b6",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"8d",x"b6",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"b6",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"4d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"ff",x"db",x"96",x"72",x"6d",x"6d",x"92",x"b6",x"b7",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b7",x"6d",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"49",x"25",x"25",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"29",x"29",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"6d",x"49",x"49",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6e",x"92",x"6e",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"6d",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"b6",x"6d",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"24",x"24",x"49",x"49",x"92",x"b6",x"6d",x"49",x"24",x"24",x"45",x"25",x"25",x"24",x"25",x"49",x"49",x"92",x"b6",x"6d",x"44",x"24",x"25",x"49",x"24",x"24",x"24",x"24",x"25",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"24",x"49",x"92",x"69",x"44",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"24",x"49",x"6d",x"92",x"6d",x"49",x"49",x"49",x"4d",x"6d",x"6e",x"b6",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"92",x"6d",x"49",x"49",x"49",x"6d",x"8e",x"b6",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"df",x"ff",x"ff",x"db",x"b6",x"b6",x"b7",x"db",x"db",x"ff",x"b6",x"91",x"6d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"db",x"db",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"b6",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"24",x"6d",x"db",x"6d",x"49",x"49",x"49",x"49",x"45",x"49"),
     (x"92",x"92",x"b6",x"db",x"ff",x"db",x"db",x"db",x"db",x"db",x"ff",x"db",x"db",x"db",x"db",x"ff",x"ff",x"db",x"92",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"92",x"49",x"49",x"49",x"69",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"92",x"ff",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"69",x"6d",x"6d",x"b6",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"8e",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"6d",x"6d",x"8d",x"d6",x"ff",x"ff",x"db",x"b6",x"b6",x"b6",x"db",x"db",x"ff",x"db",x"92",x"49",x"49",x"49",x"6d",x"6d",x"49",x"49",x"6d",x"49",x"49",x"49",x"92",x"ff",x"db",x"b6",x"92",x"92",x"6e",x"92",x"92",x"b6",x"b6",x"6e",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"b6",x"49",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"d7",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6e",x"49",x"24",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"25",x"24",x"24",x"24",x"24",x"24",x"69",x"49",x"24",x"24",x"24",x"49",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"6d",x"6e",x"92",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"24",x"24",x"20",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"8e",x"92",x"6d",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"49",x"6d",x"6d",x"92",x"6d",x"49",x"49",x"24",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"24",x"24",x"6d",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"49",x"92",x"b6",x"6d",x"45",x"24",x"45",x"45",x"49",x"6d",x"49",x"24",x"24",x"49",x"6d",x"b6",x"8e",x"49",x"49",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"24",x"6e",x"b6",x"69",x"49",x"49",x"49",x"49",x"45",x"24",x"45",x"49",x"25",x"24",x"49",x"92",x"6d",x"44",x"49",x"45",x"49",x"49",x"49",x"49",x"25",x"24",x"49",x"92",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"6e",x"b6",x"db",x"8d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"92",x"6d",x"6d",x"6d",x"6e",x"b2",x"db",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"db",x"b6",x"b6",x"92",x"b6",x"b6",x"db",x"ff",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"b6",x"ff",x"ff",x"ff",x"db",x"b6",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"8d",x"6d",x"6d",x"92",x"91",x"6d",x"6d",x"b6",x"fb",x"ff",x"db",x"6d",x"6d",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"d6",x"91",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"44",x"24",x"49",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49"),
     (x"92",x"92",x"b6",x"b6",x"db",x"ff",x"db",x"db",x"db",x"db",x"fb",x"ff",x"db",x"db",x"db",x"db",x"ff",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"ff",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"db",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b6",x"ff",x"ff",x"db",x"92",x"6d",x"69",x"69",x"6d",x"6d",x"8d",x"db",x"b6",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"92",x"49",x"49",x"49",x"49",x"69",x"69",x"6d",x"6d",x"6d",x"6d",x"92",x"d6",x"ff",x"ff",x"db",x"b6",x"92",x"b6",x"b6",x"db",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"6d",x"49",x"49",x"49",x"49",x"49",x"69",x"92",x"ff",x"df",x"b6",x"92",x"6d",x"6d",x"6d",x"6d",x"92",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"b6",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"db",x"b7",x"6e",x"6d",x"49",x"49",x"49",x"49",x"49",x"6d",x"96",x"92",x"49",x"25",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"69",x"49",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"92",x"92",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"25",x"49",x"6d",x"49",x"25",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"49",x"49",x"49",x"49",x"25",x"24",x"25",x"49",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"45",x"49",x"45",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"6d",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"20",x"00",x"20",x"24",x"24",x"24",x"24",x"24",x"00",x"20",x"24",x"24",x"24",x"49",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"00",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"92",x"6d",x"24",x"24",x"24",x"24",x"24",x"24",x"49",x"24",x"24",x"24",x"24",x"69",x"b6",x"6d",x"49",x"24",x"24",x"49",x"25",x"49",x"49",x"49",x"24",x"24",x"49",x"92",x"b6",x"49",x"49",x"49",x"45",x"24",x"24",x"25",x"24",x"24",x"24",x"24",x"92",x"b6",x"49",x"49",x"49",x"49",x"49",x"24",x"24",x"49",x"49",x"24",x"24",x"49",x"72",x"6d",x"24",x"44",x"24",x"45",x"44",x"49",x"44",x"24",x"49",x"92",x"92",x"6d",x"49",x"25",x"25",x"25",x"25",x"49",x"6d",x"b6",x"db",x"6d",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"b6",x"92",x"92",x"6e",x"92",x"92",x"b7",x"ff",x"ff",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"92",x"db",x"ff",x"db",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"49",x"49",x"49",x"49",x"6d",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"ff",x"ff",x"ff",x"b6",x"92",x"92",x"92",x"92",x"92",x"b6",x"db",x"db",x"b6",x"8d",x"8d",x"6d",x"91",x"92",x"6d",x"6d",x"b6",x"db",x"ff",x"db",x"8d",x"6d",x"6d",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"b6",x"92",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"24",x"44",x"b6",x"b6",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49")

);


begin

process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(oCoord_Y , oCoord_X);	--get from colors table 
			drawing_request	<= '1' ; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;		
		