library IEEE;
use IEEE.STD_LOGIC_1164.all;
--use IEEE.std_logic_unsigned.all;
--use ieee.numeric_std.all;
--use ieee.std_logic_arith.all;
-- Alex Grinshpun April 2017
-- Dudy Nov 13 2017


entity METRONOM_stat is
port 	(
		--////////////////////	Clock Input	 	////////////////////	
	   	CLK  		: in std_logic;
		RESETn		: in std_logic;
		oCoord_X	: in integer;
		oCoord_Y	: in integer;
		
		drawing_request	: out std_logic ;
		mVGA_RGB 	: out std_logic_vector(7 downto 0) 
	);
end METRONOM_stat;

architecture behav of METRONOM_stat is 

constant object_X_size : integer := 200;
constant object_Y_size : integer := 200;
--constant R_high		: integer := 7;
--constant R_low		: integer := 5;
--constant G_high		: integer := 4;
--constant G_low		: integer := 2;
--constant B_high		: integer := 1;
--constant B_low		: integer := 0;

type ram_array is array(0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic_vector(7 downto 0);  

-- 8 bit - color definition : "RRRGGGBB"  
constant object_colors: ram_array := ( 

(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"97",x"97",x"97",x"97",x"97",x"97",x"97",x"97",x"97",x"97",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"93",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"73",x"93",x"97",x"97",x"b7",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"bb",x"b7",x"b7",x"72",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"6e",x"72",x"97",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"bb",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"4e",x"6e",x"97",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"bb",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"72",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"bb",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2e",x"2a",x"2a",x"2a",x"4e",x"4a",x"4a",x"4e",x"2a",x"4a",x"2a",x"2a",x"2a",x"4a",x"4a",x"6e",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"db",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"2a",x"2a",x"6e",x"72",x"72",x"4e",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"2a",x"72",x"6e",x"72",x"72",x"4a",x"2a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"72",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"bb",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"49",x"92",x"92",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"72",x"49",x"92",x"72",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"db",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"4d",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"4e",x"92",x"4e",x"72",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2d",x"2d",x"4d",x"4d",x"2d",x"29",x"4d",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"92",x"6e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"52",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"4e",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"96",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"51",x"51",x"4d",x"71",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"49",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"51",x"51",x"51",x"51",x"51",x"51",x"71",x"71",x"72",x"72",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"72",x"72",x"92",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4d",x"51",x"51",x"51",x"4d",x"4d",x"71",x"71",x"71",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"51",x"51",x"51",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2e",x"2d",x"2d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4d",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2d",x"2d",x"2d",x"2d",x"2d",x"2d",x"4d",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"92",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2e",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4e",x"4a",x"4a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4a",x"4a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"4a",x"49",x"49",x"49",x"4a",x"4a",x"4a",x"4a",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"72",x"6d",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"71",x"71",x"6d",x"6d",x"6d",x"92",x"6d",x"6d",x"6d",x"92",x"92",x"91",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"25",x"25",x"25",x"29",x"29",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"49",x"49",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"92",x"71",x"6d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6d",x"72",x"92",x"92",x"92",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"6d",x"6d",x"71",x"92",x"92",x"92",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b7",x"72",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"92",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"92",x"92",x"92",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"b6",x"72",x"4e",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"92",x"92",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"49",x"b6",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"92",x"72",x"72",x"72",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"71",x"72",x"92",x"72",x"72",x"72",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"b6",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"6d",x"92",x"72",x"72",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"b6",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"72",x"72",x"6e",x"6d",x"6d",x"72",x"6e",x"72",x"72",x"72",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"72",x"72",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"92",x"72",x"72",x"92",x"72",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"52",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"49",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"6e",x"4e",x"2a",x"2a",x"4e",x"4e",x"6e",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"72",x"2a",x"2a",x"6e",x"4e",x"72",x"6e",x"6e",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"4e",x"4e",x"6e",x"4e",x"2a",x"6e",x"6e",x"92",x"72",x"6e",x"4e",x"2a",x"2a",x"6e",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"4e",x"2a",x"4e",x"6e",x"4e",x"4e",x"6e",x"29",x"72",x"92",x"92",x"92",x"6e",x"4a",x"4a",x"6e",x"92",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"96",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"72",x"4e",x"4e",x"6e",x"4e",x"4a",x"72",x"2a",x"6e",x"92",x"92",x"92",x"6e",x"4a",x"4e",x"92",x"92",x"6e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"49",x"b6",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"4e",x"4e",x"72",x"4e",x"6e",x"6e",x"6e",x"72",x"2a",x"72",x"72",x"72",x"72",x"4e",x"4e",x"72",x"92",x"92",x"92",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"b7",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"49",x"6e",x"4e",x"4e",x"6e",x"72",x"6e",x"2a",x"4e",x"4e",x"6e",x"6e",x"4e",x"4e",x"72",x"92",x"92",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"6d",x"92",x"bb",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"6e",x"72",x"4e",x"4e",x"4e",x"6e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"6e",x"92",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"b6",x"bb",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"4e",x"4e",x"6e",x"72",x"92",x"92",x"92",x"72",x"6e",x"4e",x"4e",x"4e",x"4e",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"72",x"6e",x"6e",x"6e",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"b7",x"b7",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"6e",x"92",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"92",x"4e",x"4a",x"4a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"92",x"96",x"96",x"96",x"97",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"b7",x"93",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"72",x"72",x"72",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"92",x"92",x"92",x"91",x"91",x"92",x"92",x"92",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"92",x"72",x"72",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"71",x"92",x"72",x"72",x"92",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"92",x"91",x"6d",x"71",x"6e",x"6e",x"6d",x"6d",x"6e",x"6d",x"92",x"92",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"92",x"72",x"72",x"92",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"92",x"92",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"92",x"71",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"6d",x"92",x"92",x"72",x"72",x"49",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6e",x"6e",x"6e",x"6e",x"6d",x"92",x"92",x"72",x"92",x"49",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"72",x"92",x"92",x"92",x"92",x"72",x"72",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"72",x"72",x"4e",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"72",x"6e",x"92",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"92",x"72",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6e",x"92",x"92",x"72",x"72",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"6e",x"72",x"6e",x"72",x"72",x"72",x"72",x"6e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"72",x"72",x"4a",x"2a",x"6e",x"72",x"72",x"72",x"72",x"2a",x"29",x"2a",x"4e",x"72",x"72",x"72",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"92",x"92",x"92",x"4a",x"4e",x"72",x"92",x"92",x"92",x"92",x"2a",x"2a",x"6e",x"92",x"92",x"96",x"92",x"92",x"92",x"92",x"72",x"4e",x"2a",x"4e",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"4e",x"2a",x"29",x"4e",x"72",x"92",x"92",x"96",x"96",x"92",x"92",x"92",x"92",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"96",x"92",x"4a",x"4e",x"92",x"96",x"96",x"96",x"92",x"29",x"4e",x"92",x"92",x"96",x"b6",x"b6",x"96",x"96",x"96",x"92",x"72",x"4e",x"4e",x"92",x"96",x"96",x"96",x"b6",x"96",x"96",x"96",x"96",x"92",x"6e",x"2a",x"2a",x"72",x"92",x"96",x"96",x"96",x"96",x"96",x"96",x"96",x"96",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"49",x"6e",x"92",x"96",x"96",x"92",x"72",x"29",x"72",x"92",x"92",x"96",x"96",x"96",x"92",x"96",x"96",x"96",x"92",x"4e",x"4e",x"92",x"96",x"96",x"b6",x"92",x"92",x"92",x"96",x"b6",x"96",x"6e",x"29",x"4e",x"72",x"96",x"96",x"96",x"92",x"92",x"72",x"72",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"49",x"6e",x"92",x"b6",x"b6",x"92",x"6e",x"29",x"72",x"92",x"96",x"96",x"92",x"72",x"92",x"96",x"b6",x"96",x"92",x"4e",x"4e",x"92",x"96",x"96",x"b6",x"72",x"6e",x"92",x"96",x"96",x"96",x"6e",x"29",x"4e",x"92",x"96",x"96",x"96",x"92",x"4e",x"4e",x"4e",x"4a",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"4d",x"72",x"96",x"b6",x"b6",x"92",x"4e",x"29",x"72",x"96",x"b6",x"96",x"92",x"4e",x"6e",x"96",x"b6",x"96",x"92",x"4e",x"4e",x"92",x"96",x"92",x"b6",x"72",x"6e",x"72",x"96",x"96",x"96",x"72",x"2a",x"4e",x"92",x"96",x"96",x"92",x"72",x"29",x"4a",x"4a",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"96",x"6e",x"92",x"96",x"b6",x"96",x"72",x"4a",x"29",x"72",x"96",x"b6",x"96",x"92",x"4e",x"6e",x"b6",x"b6",x"b6",x"92",x"4e",x"4e",x"92",x"b6",x"b6",x"b6",x"92",x"6e",x"92",x"b6",x"b6",x"96",x"72",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"72",x"29",x"72",x"72",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"96",x"96",x"96",x"96",x"b6",x"92",x"6e",x"2a",x"2a",x"72",x"96",x"b6",x"b6",x"92",x"4e",x"6e",x"b6",x"b6",x"b6",x"92",x"4e",x"4e",x"92",x"b6",x"b6",x"b6",x"b6",x"96",x"b6",x"b6",x"96",x"92",x"4e",x"29",x"4e",x"72",x"96",x"b6",x"96",x"72",x"49",x"92",x"96",x"96",x"96",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"96",x"96",x"96",x"96",x"92",x"92",x"4e",x"2a",x"2a",x"72",x"92",x"b6",x"b6",x"92",x"4e",x"6e",x"b6",x"96",x"b6",x"92",x"4e",x"4e",x"92",x"b6",x"92",x"b6",x"b6",x"b6",x"b6",x"96",x"92",x"6e",x"29",x"29",x"4e",x"92",x"b6",x"96",x"92",x"72",x"49",x"92",x"96",x"96",x"96",x"92",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"72",x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"96",x"92",x"96",x"96",x"b6",x"92",x"72",x"4a",x"2a",x"72",x"96",x"b6",x"b6",x"92",x"4e",x"6e",x"b6",x"b6",x"b6",x"92",x"4e",x"4e",x"92",x"96",x"96",x"b6",x"96",x"96",x"b6",x"b6",x"92",x"92",x"4e",x"29",x"4e",x"92",x"96",x"96",x"92",x"72",x"4d",x"92",x"96",x"96",x"96",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4a",x"2a",x"4e",x"72",x"6e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"96",x"92",x"6e",x"92",x"96",x"b6",x"96",x"72",x"4e",x"29",x"72",x"96",x"b6",x"96",x"92",x"4e",x"6e",x"b6",x"b6",x"b6",x"92",x"4e",x"4e",x"92",x"b6",x"b6",x"b6",x"92",x"92",x"92",x"b6",x"96",x"92",x"6e",x"29",x"4e",x"92",x"96",x"96",x"96",x"72",x"49",x"92",x"96",x"96",x"96",x"92",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"6e",x"6e",x"4a",x"4e",x"72",x"4e",x"6e",x"4e",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"29",x"4e",x"4e",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"4d",x"72",x"92",x"96",x"96",x"92",x"6e",x"29",x"72",x"96",x"96",x"96",x"92",x"4e",x"6e",x"b6",x"b6",x"96",x"92",x"4e",x"4e",x"92",x"b6",x"b6",x"96",x"72",x"72",x"92",x"96",x"b6",x"96",x"72",x"49",x"4e",x"92",x"96",x"96",x"96",x"92",x"49",x"92",x"96",x"b6",x"96",x"92",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"6e",x"72",x"4e",x"4e",x"72",x"4e",x"4e",x"6e",x"2a",x"2a",x"4e",x"4e",x"2a",x"29",x"4a",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"96",x"4d",x"6e",x"92",x"96",x"96",x"96",x"72",x"29",x"72",x"96",x"96",x"96",x"92",x"6e",x"72",x"b6",x"b6",x"96",x"92",x"4e",x"4e",x"92",x"96",x"b6",x"96",x"6e",x"6e",x"92",x"96",x"b6",x"b6",x"96",x"4e",x"4e",x"92",x"96",x"96",x"b6",x"92",x"6e",x"92",x"96",x"b6",x"96",x"92",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"29",x"6e",x"72",x"72",x"4e",x"4e",x"6e",x"4e",x"49",x"6e",x"2a",x"4e",x"4e",x"4e",x"2a",x"2a",x"72",x"72",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"b6",x"92",x"4d",x"6e",x"92",x"96",x"96",x"96",x"92",x"29",x"72",x"96",x"96",x"b6",x"96",x"92",x"92",x"b6",x"b6",x"96",x"92",x"4e",x"4e",x"92",x"96",x"b6",x"96",x"6e",x"4e",x"72",x"96",x"96",x"96",x"96",x"4e",x"4e",x"72",x"96",x"96",x"b6",x"96",x"92",x"96",x"96",x"b6",x"96",x"92",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"4e",x"2a",x"29",x"72",x"4e",x"2a",x"2a",x"4e",x"72",x"4e",x"6e",x"4e",x"6e",x"4e",x"2a",x"29",x"4e",x"72",x"72",x"72",x"4e",x"2a",x"4e",x"4e",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"96",x"96",x"4e",x"4e",x"92",x"96",x"92",x"96",x"92",x"4a",x"6e",x"96",x"96",x"96",x"96",x"96",x"96",x"b6",x"96",x"96",x"72",x"4e",x"4e",x"92",x"96",x"96",x"96",x"72",x"4e",x"6e",x"96",x"96",x"96",x"96",x"72",x"4e",x"72",x"96",x"96",x"96",x"b6",x"96",x"96",x"96",x"96",x"96",x"92",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"4e",x"72",x"92",x"6e",x"29",x"6e",x"4e",x"4a",x"2a",x"4e",x"72",x"92",x"6e",x"6e",x"4e",x"4a",x"2a",x"4e",x"72",x"4e",x"72",x"4a",x"29",x"4e",x"72",x"72",x"4e",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"96",x"96",x"92",x"4e",x"4e",x"72",x"96",x"96",x"96",x"92",x"4e",x"2a",x"72",x"92",x"96",x"96",x"96",x"96",x"96",x"96",x"92",x"4e",x"2a",x"4e",x"92",x"96",x"96",x"97",x"72",x"4a",x"4e",x"92",x"96",x"96",x"96",x"72",x"4a",x"4e",x"72",x"92",x"96",x"96",x"92",x"96",x"96",x"96",x"96",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"6e",x"6e",x"72",x"72",x"72",x"4e",x"72",x"4e",x"4a",x"4e",x"4e",x"4e",x"4e",x"6e",x"4e",x"2a",x"2a",x"4e",x"72",x"6e",x"6e",x"4a",x"6e",x"72",x"72",x"4e",x"4e",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"6e",x"6e",x"6e",x"4a",x"29",x"4e",x"6e",x"6e",x"6e",x"6e",x"4e",x"29",x"2a",x"4e",x"6e",x"72",x"72",x"72",x"72",x"4e",x"4a",x"2a",x"2a",x"2a",x"4e",x"6e",x"6e",x"6e",x"4e",x"29",x"4a",x"4e",x"6e",x"6e",x"6e",x"4e",x"2a",x"29",x"4a",x"4e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"4e",x"72",x"92",x"92",x"92",x"6e",x"72",x"6e",x"4e",x"6e",x"72",x"6e",x"4e",x"72",x"72",x"4e",x"4e",x"4e",x"4e",x"4e",x"72",x"4e",x"72",x"92",x"72",x"4e",x"2a",x"2e",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"4e",x"72",x"72",x"72",x"6e",x"6e",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"4e",x"4a",x"4a",x"4a",x"6e",x"4e",x"4e",x"4e",x"4e",x"29",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"2a",x"2a",x"29",x"29",x"2a",x"29",x"29",x"29",x"2a",x"2a",x"29",x"29",x"29",x"2a",x"29",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"2a",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"29",x"29",x"4a",x"6e",x"72",x"6e",x"4e",x"6e",x"72",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"92",x"6e",x"4a",x"2a",x"6e",x"4e",x"4a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4a",x"29",x"4a",x"4e",x"29",x"4a",x"4e",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4a",x"29",x"4a",x"4e",x"4e",x"4a",x"2a",x"2a",x"4e",x"2a",x"29",x"4e",x"4e",x"2a",x"4a",x"4e",x"4e",x"2a",x"4e",x"4e",x"4e",x"4e",x"4a",x"4e",x"4e",x"4e",x"4a",x"2a",x"2a",x"4e",x"4e",x"4e",x"29",x"2a",x"29",x"4a",x"4e",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"4e",x"4e",x"4e",x"2a",x"4e",x"4e",x"2a",x"4a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"73",x"4e",x"29",x"4a",x"2a",x"4a",x"6e",x"6e",x"4e",x"72",x"72",x"72",x"92",x"6d",x"92",x"92",x"92",x"92",x"72",x"6e",x"72",x"72",x"6e",x"2a",x"4e",x"6e",x"4e",x"4e",x"6e",x"72",x"72",x"72",x"4e",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"6e",x"29",x"72",x"72",x"4a",x"4e",x"72",x"4e",x"4e",x"72",x"72",x"4e",x"72",x"72",x"92",x"72",x"6e",x"29",x"72",x"72",x"72",x"4e",x"4e",x"6e",x"92",x"4a",x"4e",x"92",x"72",x"4e",x"6e",x"92",x"72",x"4e",x"72",x"92",x"92",x"72",x"6e",x"72",x"72",x"72",x"6e",x"4e",x"6e",x"72",x"72",x"72",x"29",x"2a",x"2a",x"6e",x"72",x"4e",x"2a",x"72",x"72",x"4a",x"4e",x"72",x"72",x"6e",x"4e",x"92",x"72",x"2a",x"6e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"6e",x"4e",x"4a",x"4e",x"6e",x"92",x"72",x"92",x"92",x"92",x"92",x"92",x"6d",x"92",x"92",x"92",x"6d",x"72",x"72",x"92",x"4a",x"29",x"4e",x"6e",x"72",x"72",x"72",x"72",x"4e",x"4e",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"96",x"92",x"49",x"92",x"92",x"49",x"6e",x"72",x"4e",x"72",x"92",x"4e",x"4a",x"72",x"72",x"72",x"72",x"72",x"49",x"92",x"6e",x"72",x"72",x"6e",x"72",x"92",x"4e",x"6e",x"92",x"72",x"4e",x"6e",x"72",x"29",x"29",x"4e",x"72",x"72",x"4e",x"4e",x"92",x"72",x"72",x"92",x"6e",x"72",x"72",x"4e",x"92",x"4e",x"2a",x"29",x"6e",x"92",x"72",x"4e",x"92",x"96",x"4a",x"72",x"72",x"4e",x"2a",x"4e",x"97",x"92",x"4a",x"6e",x"92",x"4e",x"2a",x"09",x"2a",x"4e",x"6e",x"93",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"4e",x"6e",x"72",x"6e",x"6e",x"72",x"6e",x"72",x"72",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"8e",x"8e",x"92",x"92",x"72",x"72",x"6e",x"29",x"29",x"4a",x"6e",x"72",x"6e",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"96",x"92",x"6e",x"92",x"92",x"49",x"6e",x"72",x"6e",x"72",x"72",x"29",x"29",x"6e",x"72",x"72",x"92",x"72",x"6e",x"92",x"4a",x"6e",x"72",x"72",x"92",x"92",x"72",x"72",x"92",x"72",x"6e",x"6e",x"92",x"4e",x"4a",x"2a",x"72",x"72",x"4e",x"4e",x"92",x"92",x"92",x"92",x"72",x"72",x"6e",x"49",x"72",x"6e",x"2a",x"29",x"6e",x"92",x"92",x"6e",x"92",x"96",x"4e",x"72",x"6e",x"4a",x"29",x"4e",x"97",x"96",x"6e",x"72",x"92",x"6e",x"2a",x"2a",x"2a",x"29",x"29",x"6e",x"4e",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"29",x"29",x"2a",x"4e",x"4e",x"6e",x"92",x"72",x"72",x"91",x"92",x"92",x"92",x"92",x"92",x"92",x"8e",x"8e",x"92",x"92",x"92",x"72",x"72",x"29",x"29",x"4e",x"4e",x"4a",x"29",x"2a",x"2a",x"4e",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"92",x"92",x"72",x"92",x"92",x"49",x"6e",x"72",x"6e",x"72",x"72",x"2a",x"2a",x"72",x"92",x"96",x"92",x"6e",x"72",x"92",x"4a",x"4e",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"72",x"6e",x"6e",x"92",x"72",x"4e",x"2a",x"72",x"72",x"4e",x"4a",x"92",x"96",x"92",x"6e",x"6e",x"72",x"6e",x"49",x"72",x"72",x"2a",x"29",x"6e",x"92",x"92",x"92",x"92",x"92",x"6e",x"72",x"6e",x"29",x"2a",x"4e",x"96",x"96",x"72",x"72",x"92",x"6e",x"4e",x"72",x"4e",x"2a",x"29",x"72",x"4e",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"4e",x"4e",x"4a",x"4a",x"4a",x"4e",x"72",x"72",x"92",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"4a",x"29",x"4a",x"4e",x"4e",x"4e",x"72",x"72",x"72",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"92",x"92",x"92",x"6e",x"92",x"49",x"6e",x"72",x"6e",x"72",x"72",x"29",x"2a",x"72",x"92",x"92",x"92",x"6e",x"6e",x"92",x"4a",x"6e",x"72",x"72",x"72",x"92",x"92",x"92",x"72",x"72",x"6e",x"6e",x"72",x"49",x"2a",x"29",x"72",x"72",x"4a",x"4a",x"72",x"72",x"92",x"72",x"6e",x"72",x"6e",x"4e",x"92",x"6e",x"2a",x"2a",x"6e",x"72",x"72",x"92",x"72",x"92",x"6e",x"92",x"72",x"4a",x"29",x"4e",x"92",x"72",x"92",x"72",x"72",x"6e",x"4a",x"4e",x"4e",x"2a",x"29",x"72",x"4e",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"72",x"92",x"6d",x"6d",x"6d",x"6d",x"6d",x"71",x"6d",x"92",x"92",x"92",x"92",x"92",x"92",x"72",x"72",x"4a",x"29",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"72",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"72",x"72",x"92",x"4e",x"92",x"4a",x"6e",x"72",x"4e",x"6e",x"92",x"4e",x"4e",x"72",x"72",x"72",x"72",x"72",x"4e",x"92",x"6e",x"72",x"72",x"6e",x"72",x"72",x"92",x"72",x"72",x"72",x"6e",x"6e",x"72",x"4e",x"4e",x"2a",x"72",x"72",x"4e",x"4a",x"72",x"72",x"6e",x"92",x"6e",x"72",x"72",x"6e",x"72",x"4e",x"2a",x"2a",x"6e",x"72",x"6e",x"92",x"6e",x"93",x"4e",x"72",x"72",x"6e",x"4e",x"4e",x"92",x"6e",x"92",x"6e",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"91",x"72",x"72",x"49",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"4e",x"72",x"49",x"72",x"4a",x"4e",x"6e",x"4e",x"4e",x"72",x"6e",x"4e",x"6e",x"6e",x"4e",x"6e",x"6e",x"29",x"6e",x"6e",x"72",x"4e",x"4e",x"6e",x"4e",x"6e",x"6e",x"4e",x"4e",x"4e",x"4e",x"72",x"6e",x"4e",x"2a",x"6e",x"6e",x"4a",x"2a",x"6e",x"4e",x"4e",x"6e",x"4e",x"4e",x"72",x"6e",x"6e",x"29",x"2a",x"2a",x"4e",x"4e",x"4e",x"6e",x"4a",x"72",x"4a",x"4e",x"6e",x"72",x"6e",x"4e",x"6e",x"4e",x"6e",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"4a",x"92",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"91",x"72",x"72",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"4a",x"29",x"4e",x"2a",x"2a",x"4e",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"2a",x"2a",x"4e",x"29",x"2a",x"4e",x"4e",x"2a",x"2a",x"2e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"2e",x"2a",x"2a",x"4a",x"2a",x"2a",x"4e",x"2a",x"2a",x"4a",x"2a",x"2a",x"4e",x"4e",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"92",x"92",x"72",x"6e",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"72",x"72",x"6d",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"72",x"72",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"72",x"72",x"6e",x"6d",x"6d",x"6d",x"6d",x"72",x"92",x"92",x"92",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"72",x"72",x"72",x"72",x"6e",x"6e",x"71",x"72",x"72",x"72",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"92",x"72",x"72",x"72",x"92",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"69",x"49",x"49",x"49",x"69",x"69",x"69",x"69",x"69",x"69",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"69",x"69",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"6e",x"72",x"92",x"97",x"b7",x"97",x"97",x"92",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"6e",x"93",x"b7",x"bb",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"97",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"bb",x"96",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"bb",x"db",x"db",x"db",x"fb",x"fb",x"f7",x"f7",x"f7",x"fb",x"db",x"db",x"db",x"db",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"db",x"db",x"db",x"db",x"d7",x"d6",x"d2",x"ce",x"ce",x"d2",x"d2",x"d6",x"db",x"db",x"db",x"db",x"db",x"b7",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"72",x"b7",x"db",x"db",x"d7",x"d6",x"d2",x"a9",x"84",x"84",x"84",x"84",x"89",x"d2",x"d6",x"f6",x"db",x"db",x"db",x"db",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"72",x"4e",x"6e",x"72",x"72",x"4e",x"4a",x"4e",x"29",x"4e",x"4e",x"4e",x"4e",x"4e",x"72",x"72",x"4e",x"29",x"6e",x"72",x"4e",x"4a",x"4e",x"29",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"b7",x"db",x"db",x"d7",x"d2",x"a9",x"a9",x"c9",x"ed",x"ed",x"ed",x"ed",x"cd",x"c9",x"a9",x"ce",x"d6",x"d7",x"db",x"db",x"db",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4a",x"29",x"4a",x"6e",x"4e",x"4a",x"4e",x"72",x"29",x"4e",x"72",x"72",x"4e",x"4e",x"72",x"4e",x"72",x"4e",x"6e",x"72",x"4e",x"4e",x"72",x"4a",x"6e",x"2a",x"29",x"2a",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"4e",x"92",x"d7",x"d7",x"d6",x"d2",x"89",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"ed",x"c9",x"ad",x"d6",x"d7",x"db",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"29",x"29",x"4e",x"4e",x"4a",x"6e",x"72",x"4a",x"4e",x"72",x"72",x"6e",x"6e",x"72",x"49",x"92",x"4e",x"72",x"72",x"6e",x"4e",x"6e",x"72",x"4e",x"4a",x"4e",x"6e",x"6e",x"6e",x"6e",x"6e",x"4e",x"2a",x"6e",x"97",x"d7",x"d6",x"d2",x"a9",x"c9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"c9",x"c9",x"ad",x"d6",x"d7",x"db",x"bb",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"4e",x"29",x"4e",x"4e",x"4e",x"72",x"6e",x"4e",x"6e",x"72",x"92",x"6e",x"6e",x"6e",x"29",x"72",x"4e",x"72",x"92",x"6e",x"4a",x"4e",x"92",x"4a",x"4a",x"72",x"92",x"92",x"92",x"92",x"92",x"4e",x"2a",x"72",x"b7",x"d7",x"d2",x"cd",x"a9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"cd",x"ad",x"d2",x"d6",x"db",x"db",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"4a",x"6e",x"2a",x"4e",x"4e",x"4e",x"92",x"6e",x"6e",x"6e",x"6e",x"72",x"72",x"6e",x"6e",x"29",x"72",x"4e",x"72",x"72",x"4e",x"4e",x"4e",x"93",x"2a",x"4a",x"72",x"96",x"96",x"96",x"96",x"92",x"4e",x"2a",x"72",x"b7",x"d6",x"d2",x"a9",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"d2",x"d6",x"d7",x"db",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"2a",x"4e",x"4e",x"4e",x"72",x"6e",x"72",x"6e",x"4e",x"72",x"6e",x"4e",x"72",x"4e",x"72",x"4e",x"72",x"6e",x"4e",x"4e",x"4a",x"97",x"2a",x"2a",x"4e",x"72",x"72",x"72",x"72",x"6e",x"4e",x"4a",x"92",x"b7",x"d6",x"b2",x"a9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"ad",x"d2",x"d7",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"48",x"49",x"49",x"49",x"49",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"29",x"4e",x"4e",x"4e",x"4e",x"4e",x"72",x"4e",x"4a",x"4e",x"4e",x"4e",x"6e",x"6e",x"4e",x"29",x"6e",x"72",x"4e",x"2a",x"4a",x"73",x"2a",x"2a",x"2a",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"92",x"b7",x"b6",x"ae",x"a9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"cd",x"ad",x"d2",x"d6",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"49",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"69",x"49",x"49",x"69",x"49",x"49",x"49",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"29",x"29",x"2a",x"4a",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"92",x"b7",x"d6",x"ae",x"a9",x"ee",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"ad",x"d2",x"d6",x"db",x"b7",x"72",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"92",x"b7",x"d6",x"b2",x"a9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"ad",x"d2",x"d7",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"49",x"29",x"29",x"29",x"29",x"29",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"29",x"2a",x"2a",x"25",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"b7",x"d6",x"d2",x"ad",x"cd",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"ae",x"d6",x"d7",x"db",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"2a",x"4a",x"4a",x"2a",x"4e",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4a",x"4e",x"4e",x"2a",x"4e",x"29",x"4e",x"4e",x"4e",x"6e",x"4e",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"96",x"d7",x"d6",x"ce",x"c9",x"ed",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"ed",x"cd",x"d2",x"d6",x"d7",x"b7",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"72",x"4e",x"6e",x"4e",x"4e",x"4e",x"29",x"2a",x"4e",x"4e",x"4e",x"2a",x"2a",x"2a",x"6e",x"4e",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"72",x"4e",x"6e",x"4e",x"6e",x"72",x"4e",x"72",x"29",x"72",x"4e",x"6e",x"6e",x"4e",x"6e",x"4e",x"2a",x"29",x"2a",x"29",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"b7",x"d6",x"d2",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"d2",x"d6",x"d7",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"4a",x"6e",x"4e",x"6e",x"72",x"72",x"72",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"72",x"2a",x"72",x"4e",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"72",x"6e",x"72",x"72",x"4e",x"72",x"49",x"72",x"4e",x"4e",x"4e",x"4a",x"6e",x"4e",x"2a",x"2a",x"4e",x"4e",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"b7",x"d7",x"d6",x"d2",x"cd",x"cd",x"ed",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"e9",x"ed",x"cd",x"d2",x"d6",x"d7",x"db",x"db",x"92",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"29",x"6e",x"4e",x"6e",x"92",x"92",x"72",x"2a",x"2a",x"2a",x"4e",x"4e",x"2a",x"2a",x"4e",x"4e",x"29",x"72",x"4e",x"2a",x"2a",x"2a",x"4e",x"2a",x"4e",x"92",x"72",x"92",x"72",x"6e",x"92",x"4a",x"72",x"4e",x"4e",x"4e",x"4a",x"6e",x"6e",x"2a",x"2a",x"72",x"92",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"b7",x"d7",x"d6",x"d2",x"d2",x"cd",x"ed",x"ed",x"e9",x"e9",x"e9",x"ed",x"ed",x"ce",x"d2",x"d6",x"d7",x"db",x"db",x"b7",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"29",x"6e",x"4e",x"6e",x"72",x"92",x"72",x"29",x"2a",x"2a",x"4e",x"6e",x"4e",x"4a",x"4e",x"29",x"2a",x"72",x"4e",x"2a",x"29",x"4a",x"6e",x"2a",x"4e",x"72",x"92",x"92",x"72",x"6e",x"92",x"49",x"92",x"4e",x"4e",x"4e",x"4e",x"6e",x"6e",x"4e",x"2a",x"72",x"92",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"97",x"db",x"d7",x"d7",x"d6",x"d2",x"d2",x"d2",x"ce",x"ce",x"ce",x"d2",x"d2",x"d2",x"d6",x"d7",x"db",x"db",x"b7",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"73",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"4a",x"6e",x"4e",x"4e",x"6e",x"6e",x"72",x"29",x"2a",x"2a",x"29",x"4e",x"6e",x"4e",x"4e",x"2a",x"2a",x"72",x"4e",x"2a",x"4a",x"4e",x"4e",x"29",x"4e",x"4e",x"72",x"72",x"6e",x"6e",x"92",x"49",x"72",x"4e",x"4e",x"4e",x"4e",x"4e",x"29",x"29",x"2a",x"4e",x"6e",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"b7",x"db",x"db",x"db",x"fb",x"f6",x"f6",x"f6",x"f6",x"f6",x"d6",x"f7",x"db",x"db",x"db",x"db",x"bb",x"72",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"4a",x"4e",x"4e",x"4a",x"72",x"29",x"2a",x"2a",x"4e",x"72",x"72",x"4e",x"4e",x"2a",x"2a",x"72",x"72",x"4e",x"4e",x"4e",x"29",x"2a",x"4e",x"4a",x"4e",x"6e",x"4e",x"4e",x"72",x"72",x"72",x"4a",x"4e",x"4e",x"4a",x"6e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"b7",x"db",x"db",x"db",x"db",x"fb",x"fb",x"fb",x"fb",x"db",x"db",x"db",x"db",x"db",x"b7",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4a",x"2a",x"2a",x"2a",x"2a",x"4e",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"4e",x"29",x"2a",x"2a",x"2a",x"4a",x"4a",x"4a",x"4e",x"2a",x"29",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"b7",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"db",x"b7",x"92",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"b7",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"29",x"2a",x"2a",x"29",x"29",x"2a",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"6e",x"72",x"97",x"b7",x"b7",x"b7",x"b7",x"b7",x"97",x"72",x"6e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"df",x"6e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"4e",x"4e",x"6e",x"72",x"6e",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"0a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"bb",x"72",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"97",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"72",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"97",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"b7",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"db",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"6e",x"97",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"bb",x"72",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4e",x"92",x"db",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2e",x"4e",x"6e",x"97",x"db",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"b7",x"96",x"72",x"4e",x"4e",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"2a",x"2a",x"2a",x"2a",x"2a",x"2a",x"4a",x"4a",x"4e",x"4e",x"4a",x"4a",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"4e",x"6e",x"92",x"97",x"bb",x"df",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"db",x"b7",x"96",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"72",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"92",x"93",x"93",x"93",x"93",x"93",x"93",x"92",x"92",x"92",x"92",x"92",x"92",x"97",x"97",x"b7",x"b7",x"bb",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff"),
(x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff",x"ff")
);
-- one bit mask  0 - off 1 dispaly 
type object_form is array (0 to object_Y_size - 1 , 0 to object_X_size - 1) of std_logic;
constant object : object_form := (



("00000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000"),
("00000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000"),
("00000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("00001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000"),
("00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000"),
("01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000"),
("01111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000"),
("00111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000"),
("00011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("00001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000"),
("00000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000"),
("00000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000"),
("00000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"),
("00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000")

);


signal		ObjectStartX	:  integer:=89;
signal 		ObjectStartY 	:  integer:=52;
		
signal bCoord_X : integer := 0;-- offset from start position 
signal bCoord_Y : integer := 0;

signal drawing_X : std_logic := '0';
signal drawing_Y : std_logic := '0';

--		
signal objectEndX : integer;
signal objectEndY : integer;

begin

-- Calculate object end boundaries
objectEndX	<= object_X_size+ObjectStartX;
objectEndY	<= object_Y_size+ObjectStartY;

-- Signals drawing_X[Y] are active when obects coordinates are being crossed

-- test if ooCoord is in the rectangle defined by Start and End 
	drawing_X	<= '1' when  (oCoord_X  >= ObjectStartX) and  (oCoord_X < objectEndX) else '0';
    drawing_Y	<= '1' when  (oCoord_Y  >= ObjectStartY) and  (oCoord_Y < objectEndY) else '0';

-- calculate offset from start corner 
	bCoord_X 	<= (oCoord_X - ObjectStartX) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 
	bCoord_Y 	<= (oCoord_Y - ObjectStartY) when ( drawing_X = '1' and  drawing_Y = '1'  ) else 0 ; 


process ( RESETn, CLK)

  		
   begin
	if RESETn = '0' then
	    mVGA_RGB	<=  (others => '0') ; 	
		drawing_request	<=  '0' ;

		elsif rising_edge(CLK) then
			mVGA_RGB	<=  object_colors(bCoord_Y , bCoord_X);	--get from colors table 
			drawing_request	<= object(bCoord_Y , bCoord_X) and drawing_X and drawing_Y ; -- get from mask table if inside rectangle  
	end if;

  end process;

		
end behav;		
		