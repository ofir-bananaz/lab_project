library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity ADSR_table is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  mux						: in std_logic_vector(1 downto 0);
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end ADSR_table;

architecture arch of ADSR_table is
constant array_size 			: integer := 256 ;
constant one : std_logic_vector:="01";
constant two : std_logic_vector:="10";
constant three : std_logic_vector:="11";

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal normal_table				: table_type;
signal long_table				: table_type;
signal short_table			: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;


begin 

 
  ADSR_table_proc: process(resetN, CLK)
    constant normal_table : table_type := (
	 
X"0000",
X"00FA",
X"01F4",
X"02EE",
X"03E8",
X"04E2",
X"05DC",
X"06D6",
X"07D0",
X"08CA",
X"09C4",
X"0ABE",
X"0BB8",
X"0CB2",
X"0DAC",
X"0EA6",
X"0FA0",
X"109A",
X"1194",
X"128E",
X"1388",
X"1482",
X"157C",
X"1676",
X"1770",
X"186A",
X"1964",
X"1A5E",
X"1B58",
X"1C52",
X"1D4C",
X"1E46",
X"1F40",
X"203A",
X"2134",
X"222E",
X"2328",
X"2422",
X"251C",
X"2616",
X"2710",
X"280A",
X"2904",
X"29FE",
X"2AF8",
X"2BF2",
X"2CEC",
X"2DE6",
X"2EE0",
X"2FDA",
X"30D4",
X"31CE",
X"32C8",
X"33C2",
X"34BC",
X"35B6",
X"36B0",
X"37AA",
X"38A4",
X"399E",
X"3A98",
X"3B92",
X"3C8C",
X"3D86",
X"3E80",
X"3E80",
X"3DCE",
X"3D1C",
X"3C6A",
X"3BB8",
X"3B07",
X"3A55",
X"39A3",
X"38F1",
X"3840",
X"378E",
X"36DC",
X"362A",
X"3578",
X"34C7",
X"3415",
X"3363",
X"32B1",
X"3200",
X"314E",
X"309C",
X"2FEA",
X"2F38",
X"2E87",
X"2DD5",
X"2D23",
X"2C71",
X"2BC0",
X"2B0E",
X"2A5C",
X"29AA",
X"28F8",
X"2847",
X"2795",
X"26E3",
X"2631",
X"2580",
X"24CE",
X"241C",
X"236A",
X"22B8",
X"2207",
X"2155",
X"20A3",
X"1FF1",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"1F40",
X"3E80",
X"3A46",
X"3655",
X"32A9",
X"2F3C",
X"2C0B",
X"2910",
X"264A",
X"23B3",
X"2149",
X"1F09",
X"1CF0",
X"1AFB",
X"1928",
X"1774",
X"15DF",
X"1464",
X"1303",
X"11BA",
X"1087",
X"0F69",
X"0E5E",
X"0D66",
X"0C7E",
X"0BA5",
X"0ADC",
X"0A20",
X"0971",
X"08CD",
X"0835",
X"07A7",
X"0722",
X"06A7",
X"0634",
X"05C8",
X"0564",
X"0507",
X"04B0",
X"045F",
X"0413",
X"03CC",
X"038B",
X"034D",
X"0314",
X"02DF",
X"02AD",
X"027F",
X"0254",
X"022B",
X"0206",
X"01E3",
X"01C2",
X"01A4",
X"0187",
X"016D",
X"0154",
X"013D",
X"0127",
X"0113",
X"0101",
X"00EF",
X"00DF",
X"00D0",
X"00C2",
X"00B5",
X"00A9",
X"009D",
X"0092",
X"0089",
X"007F",
X"0077",
X"006F",
X"0067",
X"0060",
X"005A",
X"0053",
X"004E",
X"0048",
X"0044",
X"003F",
X"003B",
X"0037",
X"0033",
X"002F",
X"002C",
X"0029",
X"0026",
X"0024",
X"0021",
X"001F",
X"001D",
X"001B",
X"0019",
X"0017",
X"0016",
X"0014",
X"0013",
X"0011",
X"0010",
X"000F",
X"000E",
X"000D",
X"000C",
X"000B",
X"000B",
X"000A",
X"0009",
X"0008"
);


constant long_table : table_type := (

X"0000",
X"0122",
X"0245",
X"0368",
X"048B",
X"05AE",
X"06D1",
X"07F4",
X"0917",
X"0A3A",
X"0B5D",
X"0C7F",
X"0DA2",
X"0EC5",
X"0FE8",
X"110B",
X"122E",
X"1351",
X"1474",
X"1597",
X"16BA",
X"17DD",
X"18FF",
X"1A22",
X"1B45",
X"1C68",
X"1D8B",
X"1EAE",
X"1FD1",
X"20F4",
X"2217",
X"233A",
X"245D",
X"2580",
X"26A2",
X"27C5",
X"28E8",
X"2A0B",
X"2B2E",
X"2C51",
X"2D74",
X"2E97",
X"2FBA",
X"30DD",
X"31FF",
X"3322",
X"3445",
X"3568",
X"368B",
X"37AE",
X"38D1",
X"39F4",
X"3B17",
X"3C3A",
X"3D5D",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3A46",
X"3655",
X"32A9",
X"2F3C",
X"2C0B",
X"2910",
X"264A",
X"23B3",
X"2149",
X"1F09",
X"1CF0",
X"1AFB",
X"1928",
X"1774",
X"15DF",
X"1464",
X"1303",
X"11BA",
X"1087",
X"0F69",
X"0E5E",
X"0D66",
X"0C7E",
X"0BA5",
X"0ADC",
X"0A20",
X"0971",
X"08CD",
X"0835",
X"07A7",
X"0722",
X"06A7",
X"0634",
X"05C8",
X"0564",
X"0507",
X"04B0",
X"045F",
X"0413",
X"03CC",
X"038B",
X"034D",
X"0314",
X"02DF",
X"02AD",
X"027F",
X"0254",
X"022B",
X"0206",
X"01E3",
X"01C2",
X"01A4",
X"0187",
X"016D",
X"0154",
X"013D",
X"0127",
X"0113",
X"0101",
X"00EF",
X"00DF",
X"00D0",
X"00C2",
X"00B5",
X"00A9",
X"009D",
X"0092",
X"0089",
X"007F",
X"0077",
X"006F",
X"0067",
X"0060",
X"005A",
X"0053",
X"004E",
X"0048",
X"0044",
X"003F",
X"003B",
X"0037",
X"0033",
X"002F",
X"002C",
X"0029",
X"0026",
X"0024",
X"0021",
X"001F",
X"001D",
X"001B",
X"0019",
X"0017",
X"0016",
X"0014",
X"0013",
X"0011",
X"0010",
X"000F",
X"000E",
X"000D",
X"000C",
X"000B",
X"000B",
X"000A",
X"0009",
X"0008",
X"0008",
X"0007",
X"0007",
X"0006",
X"0006",
X"0005",
X"0005",
X"0005",
X"0004",
X"0004",
X"0004",
X"0003",
X"0003",
X"0003",
X"0003",
X"0002",
X"0002",
X"0002",
X"0002",
X"0002",
X"0002",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0001",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000");

constant short_table : table_type := (

X"0000",
X"00A0",
X"0140",
X"01E0",
X"0280",
X"0320",
X"03C0",
X"0460",
X"0500",
X"05A0",
X"0640",
X"06E0",
X"0780",
X"0820",
X"08C0",
X"0960",
X"0A00",
X"0AA0",
X"0B40",
X"0BE0",
X"0C80",
X"0D20",
X"0DC0",
X"0E60",
X"0F00",
X"0FA0",
X"1040",
X"10E0",
X"1180",
X"1220",
X"12C0",
X"1360",
X"1400",
X"14A0",
X"1540",
X"15E0",
X"1680",
X"1720",
X"17C0",
X"1860",
X"1900",
X"19A0",
X"1A40",
X"1AE0",
X"1B80",
X"1C20",
X"1CC0",
X"1D60",
X"1E00",
X"1EA0",
X"1F40",
X"1FE0",
X"2080",
X"2120",
X"21C0",
X"2260",
X"2300",
X"23A0",
X"2440",
X"24E0",
X"2580",
X"2620",
X"26C0",
X"2760",
X"2800",
X"28A0",
X"2940",
X"29E0",
X"2A80",
X"2B20",
X"2BC0",
X"2C60",
X"2D00",
X"2DA0",
X"2E40",
X"2EE0",
X"2F80",
X"3020",
X"30C0",
X"3160",
X"3200",
X"32A0",
X"3340",
X"33E0",
X"3480",
X"3520",
X"35C0",
X"3660",
X"3700",
X"37A0",
X"3840",
X"38E0",
X"3980",
X"3A20",
X"3AC0",
X"3B60",
X"3C00",
X"3CA0",
X"3D40",
X"3DE0",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"47E4",
X"4308",
X"3E80",
X"3A46",
X"3655",
X"32A9",
X"2F3C",
X"2C0B",
X"2910",
X"264A",
X"23B3",
X"2149",
X"1F09",
X"1CF0",
X"1AFB",
X"1928",
X"1774",
X"15DF",
X"1464",
X"1303",
X"11BA",
X"1087",
X"0F69",
X"0E5E",
X"0D66",
X"0C7E",
X"0BA5",
X"0ADC",
X"0A20",
X"0971",
X"08CD",
X"0835",
X"07A7",
X"0722",
X"06A7",
X"0634",
X"05C8",
X"0564",
X"0507",
X"04B0",
X"045F",
X"0413",
X"03CC",
X"038B",
X"034D",
X"0314",
X"02DF",
X"02AD",
X"027F",
X"0254",
X"022B",
X"0206",
X"01E3",
X"01C2",
X"01A4",
X"0187",
X"016D",
X"0154",
X"013D",
X"0127",
X"0113",
X"0101",
X"00EF",
X"00DF",
X"00D0",
X"00C2",
X"00B5",
X"00A9",
X"009D",
X"0092",
X"0089",
X"007F",
X"0077",
X"006F",
X"0067",
X"0060",
X"005A",
X"0053",
X"004E",
X"0048",
X"0044",
X"003F",
X"003B",
X"0037",
X"0033",
X"002F",
X"002C",
X"0029",
X"0026",
X"0024",
X"0021",
X"001F",
X"001D",
X"001B",
X"0019",
X"0017",
X"0016",
X"0014",
X"0013",
X"0011",
X"0010",
X"000F",
X"000E",
X"000D",
X"000C",
X"000B",
X"000B",
X"000A",
X"0009",
X"0008",
X"0008",
X"0007",
X"0007",
X"0006",
X"0006",
X"0005",
X"0005",
X"0005",
X"0004",
X"0004",
X"0004",
X"0003",
X"0003",
X"0003",
X"0003",
X"0002",
X"0002",
X"0002",
X"0002");

begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
    elsif(rising_edge(CLK)) then
		case mux is
			when two =>
				Q_tmp <= short_table(conv_integer(ADDR));
			when three => 
				Q_tmp <= long_table(conv_integer(ADDR));
			when others=>
				Q_tmp <= normal_table(conv_integer(ADDR));
		end case;
   end if;
  end process;
 Q <= Q_tmp; 
		   
end arch;
