--------------------------------------
-- SinTable.vhd
-- Written by Gadi and Eran Tuchman.
-- All rights reserved, Copyright 2009
--------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;

entity sintable is
port(
  CLK     					: in std_logic;
  resetN 					: in std_logic;
  wave						: in std_logic_vector(2 downto 0);
  ADDR    					: in std_logic_vector(7 downto 0);
  Q       					: out std_logic_vector(15 downto 0)
);
end sintable;

architecture arch of sintable is
constant array_size 			: integer := 256 ;
constant ZERO : std_logic_vector:="000";
constant one : std_logic_vector:="001";
constant two : std_logic_vector:="010";
constant three : std_logic_vector:="100";

type table_type is array(0 to array_size - 1) of std_logic_vector(15 downto 0);
signal sin_table				: table_type;
signal sincos_table				: table_type;
signal square_table			: table_type;
signal Q_tmp       			:  std_logic_vector(15 downto 0) ;
SIGNAL COMP 					:	STD_LOGIC_VECTOR(2 DOWNTO 0);

begin
 
   
  sintable_proc: process(resetN, CLK)
    constant sin_table : table_type := (
---start 0 v
X"0000",
X"0188",
X"0311",
X"0499",
X"0620",
X"07A6",
X"092B",
X"0AAF",
X"0C31",
X"0DB1",
X"0F2F",
X"10AB",
X"1224",
X"139A",
X"150E",
X"167E",
X"17EA",
X"1953",
X"1AB8",
X"1C19",
X"1D76",
X"1ECE",
X"2021",
X"216F",
X"22B9",
X"23FC",
X"253B",
X"2673",
X"27A6",
X"28D2",
X"29F8",
X"2B18",
X"2C31",
X"2D43",
X"2E4F",
X"2F53",
X"3050",
X"3145",
X"3233",
X"3319",
X"33F7",
X"34CD",
X"359B",
X"3661",
X"371E",
X"37D3",
X"387F",
X"3923",
X"39BE",
X"3A4F",
X"3AD8",
X"3B58",
X"3BCF",
X"3C3C",
X"3CA0",
X"3CFB",
X"3D4C",
X"3D94",
X"3DD2",
X"3E07",
X"3E32",
X"3E54",
X"3E6C",
X"3E7B",
X"3E80",
X"3E7B",
X"3E6C",
X"3E54",
X"3E32",
X"3E07",
X"3DD2",
X"3D94",
X"3D4C",
X"3CFB",
X"3CA0",
X"3C3C",
X"3BCF",
X"3B58",
X"3AD8",
X"3A4F",
X"39BE",
X"3923",
X"387F",
X"37D3",
X"371E",
X"3661",
X"359B",
X"34CD",
X"33F7",
X"3319",
X"3233",
X"3145",
X"3050",
X"2F53",
X"2E4F",
X"2D43",
X"2C31",
X"2B18",
X"29F8",
X"28D2",
X"27A6",
X"2673",
X"253B",
X"23FC",
X"22B9",
X"216F",
X"2021",
X"1ECE",
X"1D76",
X"1C19",
X"1AB8",
X"1953",
X"17EA",
X"167E",
X"150E",
X"139A",
X"1224",
X"10AB",
X"0F2F",
X"0DB1",
X"0C31",
X"0AAF",
X"092B",
X"07A6",
X"0620",
X"0499",
X"0311",
X"0188",
X"0000",
X"FE78",
X"FCEF",
X"FB67",
X"F9E0",
X"F85A",
X"F6D5",
X"F551",
X"F3CF",
X"F24F",
X"F0D1",
X"EF55",
X"EDDC",
X"EC66",
X"EAF2",
X"E982",
X"E816",
X"E6AD",
X"E548",
X"E3E7",
X"E28A",
X"E132",
X"DFDF",
X"DE91",
X"DD47",
X"DC04",
X"DAC5",
X"D98D",
X"D85A",
X"D72E",
X"D608",
X"D4E8",
X"D3CF",
X"D2BD",
X"D1B1",
X"D0AD",
X"CFB0",
X"CEBB",
X"CDCD",
X"CCE7",
X"CC09",
X"CB33",
X"CA65",
X"C99F",
X"C8E2",
X"C82D",
X"C781",
X"C6DD",
X"C642",
X"C5B1",
X"C528",
X"C4A8",
X"C431",
X"C3C4",
X"C360",
X"C305",
X"C2B4",
X"C26C",
X"C22E",
X"C1F9",
X"C1CE",
X"C1AC",
X"C194",
X"C185",
X"C180",
X"C185",
X"C194",
X"C1AC",
X"C1CE",
X"C1F9",
X"C22E",
X"C26C",
X"C2B4",
X"C305",
X"C360",
X"C3C4",
X"C431",
X"C4A8",
X"C528",
X"C5B1",
X"C642",
X"C6DD",
X"C781",
X"C82D",
X"C8E2",
X"C99F",
X"CA65",
X"CB33",
X"CC09",
X"CCE7",
X"CDCD",
X"CEBB",
X"CFB0",
X"D0AD",
X"D1B1",
X"D2BD",
X"D3CF",
X"D4E8",
X"D608",
X"D72E",
X"D85A",
X"D98D",
X"DAC5",
X"DC04",
X"DD47",
X"DE91",
X"DFDF",
X"E132",
X"E28A",
X"E3E7",
X"E548",
X"E6AD",
X"E816",
X"E982",
X"EAF2",
X"EC66",
X"EDDC",
X"EF55",
X"F0D1",
X"F24F",
X"F3CF",
X"F551",
X"F6D5",
X"F85A",
X"F9E0",
X"FB67",
X"FCEF",
X"FE78"
 );
 

    constant sincos_table : table_type := (
X"0000",
X"0310",
X"061E",
X"0925",
X"0C22",
X"0F12",
X"11F2",
X"14BE",
X"1775",
X"1A12",
X"1C94",
X"1EF7",
X"213A",
X"235A",
X"2554",
X"2728",
X"28D4",
X"2A56",
X"2BAC",
X"2CD7",
X"2DD4",
X"2EA4",
X"2F47",
X"2FBB",
X"3002",
X"301C",
X"3009",
X"2FCB",
X"2F62",
X"2ED0",
X"2E16",
X"2D35",
X"2C31",
X"2B0B",
X"29C5",
X"2861",
X"26E3",
X"254C",
X"23A0",
X"21E2",
X"2014",
X"1E3A",
X"1C56",
X"1A6C",
X"187F",
X"1692",
X"14A8",
X"12C4",
X"10E9",
X"0F1B",
X"0D5B",
X"0BAD",
X"0A14",
X"0891",
X"0728",
X"05DA",
X"04AA",
X"0399",
X"02A9",
X"01DB",
X"0131",
X"00AC",
X"004C",
X"0013",
X"0000",
X"0013",
X"004C",
X"00AC",
X"0131",
X"01DB",
X"02A9",
X"0399",
X"04AA",
X"05DA",
X"0728",
X"0891",
X"0A14",
X"0BAD",
X"0D5B",
X"0F1B",
X"10E9",
X"12C4",
X"14A8",
X"1692",
X"187F",
X"1A6C",
X"1C56",
X"1E3A",
X"2014",
X"21E2",
X"23A0",
X"254C",
X"26E3",
X"2861",
X"29C5",
X"2B0B",
X"2C31",
X"2D35",
X"2E16",
X"2ED0",
X"2F62",
X"2FCB",
X"3009",
X"301C",
X"3002",
X"2FBB",
X"2F47",
X"2EA4",
X"2DD4",
X"2CD7",
X"2BAC",
X"2A56",
X"28D4",
X"2728",
X"2554",
X"235A",
X"213A",
X"1EF7",
X"1C94",
X"1A12",
X"1775",
X"14BE",
X"11F2",
X"0F12",
X"0C22",
X"0925",
X"061E",
X"0310",
X"0000",
X"FCF0",
X"F9E2",
X"F6DB",
X"F3DE",
X"F0EE",
X"EE0E",
X"EB42",
X"E88B",
X"E5EE",
X"E36C",
X"E109",
X"DEC6",
X"DCA6",
X"DAAC",
X"D8D8",
X"D72C",
X"D5AA",
X"D454",
X"D329",
X"D22C",
X"D15C",
X"D0B9",
X"D045",
X"CFFE",
X"CFE4",
X"CFF7",
X"D035",
X"D09E",
X"D130",
X"D1EA",
X"D2CB",
X"D3CF",
X"D4F5",
X"D63B",
X"D79F",
X"D91D",
X"DAB4",
X"DC60",
X"DE1E",
X"DFEC",
X"E1C6",
X"E3AA",
X"E594",
X"E781",
X"E96E",
X"EB58",
X"ED3C",
X"EF17",
X"F0E5",
X"F2A5",
X"F453",
X"F5EC",
X"F76F",
X"F8D8",
X"FA26",
X"FB56",
X"FC67",
X"FD57",
X"FE25",
X"FECF",
X"FF54",
X"FFB4",
X"FFED",
X"0000",
X"FFED",
X"FFB4",
X"FF54",
X"FECF",
X"FE25",
X"FD57",
X"FC67",
X"FB56",
X"FA26",
X"F8D8",
X"F76F",
X"F5EC",
X"F453",
X"F2A5",
X"F0E5",
X"EF17",
X"ED3C",
X"EB58",
X"E96E",
X"E781",
X"E594",
X"E3AA",
X"E1C6",
X"DFEC",
X"DE1E",
X"DC60",
X"DAB4",
X"D91D",
X"D79F",
X"D63B",
X"D4F5",
X"D3CF",
X"D2CB",
X"D1EA",
X"D130",
X"D09E",
X"D035",
X"CFF7",
X"CFE4",
X"CFFE",
X"D045",
X"D0B9",
X"D15C",
X"D22C",
X"D329",
X"D454",
X"D5AA",
X"D72C",
X"D8D8",
X"DAAC",
X"DCA6",
X"DEC6",
X"E109",
X"E36C",
X"E5EE",
X"E88B",
X"EB42",
X"EE0E",
X"F0EE",
X"F3DE",
X"F6DB",
X"F9E2",
X"FCF0");


    constant square_table : table_type := (
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"0000",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80",
X"3E80");

 
 begin

    if (resetN='0') then
		Q_tmp <= ( others => '0');
		COMP<= ZERO;
    elsif(rising_edge(CLK)) then
		IF(COMP/=WAVE AND WAVE/=ZERO) THEN
			COMP<=WAVE;
		END IF;
		
		CASE COMP IS
			WHEN TWO =>
					Q_tmp <= sincos_table(conv_integer(ADDR));
			when three => 
				Q_tmp <= square_table(conv_integer(ADDR));
			when others=>
				Q_tmp <= sin_table(conv_integer(ADDR));
		END CASE;
   end if;
  end process;
 Q <= Q_tmp; 
		   
end arch;